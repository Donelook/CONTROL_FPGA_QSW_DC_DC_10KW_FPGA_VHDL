-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 25 2024 17:56:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    error_pin : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__53311\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53309\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53291\ : std_logic;
signal \N__53290\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53281\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53273\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53263\ : std_logic;
signal \N__53262\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53246\ : std_logic;
signal \N__53245\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53236\ : std_logic;
signal \N__53235\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53227\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53210\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53208\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53182\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53172\ : std_logic;
signal \N__53169\ : std_logic;
signal \N__53168\ : std_logic;
signal \N__53163\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53146\ : std_logic;
signal \N__53143\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53134\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53112\ : std_logic;
signal \N__53111\ : std_logic;
signal \N__53108\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53073\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53062\ : std_logic;
signal \N__53059\ : std_logic;
signal \N__53056\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53023\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52977\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52968\ : std_logic;
signal \N__52965\ : std_logic;
signal \N__52962\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52945\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52938\ : std_logic;
signal \N__52935\ : std_logic;
signal \N__52932\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52921\ : std_logic;
signal \N__52920\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52918\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52865\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52855\ : std_logic;
signal \N__52852\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52834\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52829\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52823\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52802\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52767\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52761\ : std_logic;
signal \N__52758\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52732\ : std_logic;
signal \N__52729\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52718\ : std_logic;
signal \N__52715\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52702\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52692\ : std_logic;
signal \N__52687\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52657\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52655\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52652\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52648\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52645\ : std_logic;
signal \N__52644\ : std_logic;
signal \N__52643\ : std_logic;
signal \N__52642\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52639\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52636\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52633\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52630\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52627\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52622\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52617\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52614\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52611\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52608\ : std_logic;
signal \N__52607\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52604\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52601\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52595\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52592\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52589\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52584\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52582\ : std_logic;
signal \N__52581\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52579\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52575\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52569\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52566\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52557\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52554\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52551\ : std_logic;
signal \N__52550\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52292\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52271\ : std_logic;
signal \N__52270\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52262\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52256\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52252\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52250\ : std_logic;
signal \N__52249\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52238\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52235\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52219\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52209\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52193\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52181\ : std_logic;
signal \N__52180\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52175\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52172\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52169\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51949\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51936\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51925\ : std_logic;
signal \N__51922\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51897\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51884\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51850\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51848\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51845\ : std_logic;
signal \N__51844\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51799\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51745\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51736\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51698\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51650\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51647\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51644\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51635\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51608\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51605\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51590\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51584\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51511\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51417\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51413\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51376\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51373\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51370\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51357\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51345\ : std_logic;
signal \N__51344\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51341\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51311\ : std_logic;
signal \N__51308\ : std_logic;
signal \N__51305\ : std_logic;
signal \N__51302\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51274\ : std_logic;
signal \N__51271\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51103\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51091\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51077\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51067\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51061\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50998\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50745\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50677\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50635\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50093\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50090\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50083\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50075\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49376\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49006\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41389\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \pwm_generator_inst.O_0_1\ : std_logic;
signal \pwm_generator_inst.O_0_0\ : std_logic;
signal \pwm_generator_inst.O_0_5\ : std_logic;
signal \pwm_generator_inst.O_0_3\ : std_logic;
signal \pwm_generator_inst.O_0_4\ : std_logic;
signal \pwm_generator_inst.O_0_2\ : std_logic;
signal \pwm_generator_inst.O_0_6\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_0\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_8\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.O_11\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_11\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_15\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_19\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_20\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_21\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_22\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_23\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_24\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_cry_25\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_19\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_21\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_22\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_23\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_25\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_20\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_24\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_15\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un18_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_8\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_15\ : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_1_26\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_\ : std_logic;
signal \pwm_generator_inst.un5_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_axb_16\ : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal \pwm_generator_inst.O_0_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_0_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_0_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.O_0_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.O_0_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.O_0_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.O_0_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0\ : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7\ : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_19\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_20\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_21\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_22\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_23\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_24\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_7\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_25\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un18_threshold1_18\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\ : std_logic;
signal \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\ : std_logic;
signal \pwm_generator_inst.N_179_i\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \pwm_generator_inst.N_180_i\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.N_181_i\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.N_182_i\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.N_183_i\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.N_184_i\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.N_185_i\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.N_186_i\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.N_187_i\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \pwm_generator_inst.N_188_i\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_0\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_8\ : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_30\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_lt28\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_16 : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_17 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_18 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_19 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_21 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_0\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_8\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_16\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_24\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counter_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0_g\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_8\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_24 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_25 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_26 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_27 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal s3_phy_c : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_ns_0_0_1_cascade_\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_1 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_6 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_5 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_13 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_7 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_4 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_2 : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_3 : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_0\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_8\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt16\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_30\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_0\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_8\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_15\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_30\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_0\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_8\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_15\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_23\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_i_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counter_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_0\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_16\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_24\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_i_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counter_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0_g\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt20\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_20 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt22\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_22 : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_23 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_i_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un6_running_lt30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\ : std_logic;
signal \phase_controller_inst2.start_flagZ0\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_4\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.state_ns_0_0_1_cascade_\ : std_logic;
signal \phase_controller_inst1.start_flagZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_14 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_12 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_11 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_8 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt28\ : std_logic;
signal phase_controller_inst1_stoper_tr_target_ticks_1_i_28 : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.counterZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un6_running_lt30\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_start_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \bfn_12_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \GB_BUFFER_reset_c_g_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_7\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_15\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_23\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_168_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_167_i\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_i_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_0\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_8\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_15\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counter\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.counterZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.control_input_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_1 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_3 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_4 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_5 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_6 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_7 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_8 : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_9 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_10 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_11 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_12 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_13 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_14 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_16 : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_17 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_18 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_19 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_20 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_21 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_22 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_23 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_24 : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_25 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_26 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_27 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_15 : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\ : std_logic;
signal phase_controller_inst1_stoper_hc_target_ticks_1_i_28 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.N_1379_i\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_165_i\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i_g\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_18_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_166_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.timer_s1.N_164_i\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal s1_phy_c : std_logic;
signal state_3 : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_145\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \pwm_generator_inst.un3_threshold_iZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_10 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_162\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_160\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal reset_c_g : std_logic;

signal reset_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    pwm_output <= pwm_output_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__37882\&\N__37855\&\N__38182\&\N__37822\&\N__37795\&\N__38209\&\N__37504\&\N__37969\&\N__38008\&\N__37912\&\N__37939\&\N__37276\&\N__37531\&\N__37306\&\N__37333\&\N__37357\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__51644\&'0'&\N__51643\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_A_wire\ <= '0'&\N__51797\&\N__51800\&\N__51798\&\N__51801\&\N__51799\&\N__51868\&\N__52663\&\N__53020\&\N__51676\&\N__53146\&\N__53062\&\N__52927\&\N__51727\&\N__51751\&\N__52990\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__51621\&'0'&\N__51620\;
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(15);
    \pwm_generator_inst.O_0_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(14);
    \pwm_generator_inst.O_0_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(13);
    \pwm_generator_inst.O_0_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(12);
    \pwm_generator_inst.O_0_11\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(11);
    \pwm_generator_inst.O_0_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(10);
    \pwm_generator_inst.O_0_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(9);
    \pwm_generator_inst.O_0_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(8);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(7);
    \pwm_generator_inst.O_0_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(6);
    \pwm_generator_inst.O_0_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(5);
    \pwm_generator_inst.O_0_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(4);
    \pwm_generator_inst.O_0_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(3);
    \pwm_generator_inst.O_0_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(2);
    \pwm_generator_inst.O_0_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(1);
    \pwm_generator_inst.O_0_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_A_wire\ <= '0'&\N__22822\&\N__22861\&\N__22897\&\N__51922\&\N__21625\&\N__21718\&\N__21673\&\N__21694\&\N__21646\&\N__21760\&\N__21739\&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&\N__51356\&\N__51372\&\N__51359\&\N__51371\&\N__51357\&'0'&'0'&\N__51370\&\N__51358\&\N__51369\;
    \pwm_generator_inst.un5_threshold_1_26\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(26);
    \pwm_generator_inst.un5_threshold_1_25\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(25);
    \pwm_generator_inst.un5_threshold_1_24\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(24);
    \pwm_generator_inst.un5_threshold_1_23\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(23);
    \pwm_generator_inst.un5_threshold_1_22\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(22);
    \pwm_generator_inst.un5_threshold_1_21\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(21);
    \pwm_generator_inst.un5_threshold_1_20\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(20);
    \pwm_generator_inst.un5_threshold_1_19\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(19);
    \pwm_generator_inst.un5_threshold_1_18\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(18);
    \pwm_generator_inst.un5_threshold_1_17\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(17);
    \pwm_generator_inst.un5_threshold_1_16\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(16);
    \pwm_generator_inst.un5_threshold_1_15\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(12);
    \pwm_generator_inst.O_11\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_A_wire\ <= \N__51851\&\N__51859\&\N__51850\&\N__51858\&\N__51849\&\N__51857\&\N__51848\&\N__51856\&\N__51847\&\N__51854\&\N__51846\&\N__51855\&\N__51845\&\N__51853\&\N__51844\&\N__51852\;
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__51170\&'0'&\N__51169\;
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\(0);
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_A_wire\ <= '0'&\N__23131\&\N__23140\&\N__23152\&\N__22927\&\N__22936\&\N__22945\&\N__22954\&\N__22963\&\N__22972\&\N__22981\&\N__22990\&\N__22687\&\N__22717\&\N__22750\&\N__22786\;
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&\N__51076\&\N__51080\&\N__51086\&\N__51079\&\N__51084\&'0'&'0'&\N__51078\&\N__51085\&\N__51077\;
    \pwm_generator_inst.un5_threshold_2_1_16\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(16);
    \pwm_generator_inst.un5_threshold_2_1_15\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(15);
    \pwm_generator_inst.un5_threshold_2_14\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(14);
    \pwm_generator_inst.un5_threshold_2_13\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(13);
    \pwm_generator_inst.un5_threshold_2_12\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(12);
    \pwm_generator_inst.un5_threshold_2_11\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(11);
    \pwm_generator_inst.un5_threshold_2_10\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(10);
    \pwm_generator_inst.un5_threshold_2_9\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(9);
    \pwm_generator_inst.un5_threshold_2_8\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(8);
    \pwm_generator_inst.un5_threshold_2_7\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(7);
    \pwm_generator_inst.un5_threshold_2_6\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(6);
    \pwm_generator_inst.un5_threshold_2_5\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(5);
    \pwm_generator_inst.un5_threshold_2_4\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(4);
    \pwm_generator_inst.un5_threshold_2_3\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(3);
    \pwm_generator_inst.un5_threshold_2_2\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(2);
    \pwm_generator_inst.un5_threshold_2_1\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(1);
    \pwm_generator_inst.un5_threshold_2_0\ <= \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__37387\&\N__37417\&\N__37444\&\N__37051\&\N__37078\&\N__37102\&\N__37129\&\N__37162\&\N__37189\&\N__37216\&\N__37243\&\N__36967\&\N__36991\&\N__37018\&\N__50218\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__51579\&'0'&\N__51578\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__24919\,
            RESETB => \N__35719\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__51645\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__51642\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__51622\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__51619\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__51360\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__51355\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_A_wire\,
            C => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_C_wire\,
            B => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__51171\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__51168\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0_O_wire\
        );

    \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__51090\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__51075\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_A_wire\,
            C => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_C_wire\,
            B => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__51494\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__51577\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__53309\,
            GLOBALBUFFEROUTPUT => reset_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53311\,
            DIN => \N__53310\,
            DOUT => \N__53309\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53311\,
            PADOUT => \N__53310\,
            PADIN => \N__53309\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53300\,
            DIN => \N__53299\,
            DOUT => \N__53298\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53300\,
            PADOUT => \N__53299\,
            PADIN => \N__53298\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53291\,
            DIN => \N__53290\,
            DOUT => \N__53289\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53291\,
            PADOUT => \N__53290\,
            PADIN => \N__53289\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53282\,
            DIN => \N__53281\,
            DOUT => \N__53280\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53282\,
            PADOUT => \N__53281\,
            PADIN => \N__53280\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__50368\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53273\,
            DIN => \N__53272\,
            DOUT => \N__53271\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53273\,
            PADOUT => \N__53272\,
            PADIN => \N__53271\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53264\,
            DIN => \N__53263\,
            DOUT => \N__53262\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53264\,
            PADOUT => \N__53263\,
            PADIN => \N__53262\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53255\,
            DIN => \N__53254\,
            DOUT => \N__53253\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53255\,
            PADOUT => \N__53254\,
            PADIN => \N__53253\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53246\,
            DIN => \N__53245\,
            DOUT => \N__53244\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53246\,
            PADOUT => \N__53245\,
            PADIN => \N__53244\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53237\,
            DIN => \N__53236\,
            DOUT => \N__53235\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53237\,
            PADOUT => \N__53236\,
            PADIN => \N__53235\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53228\,
            DIN => \N__53227\,
            DOUT => \N__53226\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53228\,
            PADOUT => \N__53227\,
            PADIN => \N__53226\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53219\,
            DIN => \N__53218\,
            DOUT => \N__53217\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53219\,
            PADOUT => \N__53218\,
            PADIN => \N__53217\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38071\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53210\,
            DIN => \N__53209\,
            DOUT => \N__53208\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53210\,
            PADOUT => \N__53209\,
            PADIN => \N__53208\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53201\,
            DIN => \N__53200\,
            DOUT => \N__53199\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53201\,
            PADOUT => \N__53200\,
            PADIN => \N__53199\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12303\ : CascadeMux
    port map (
            O => \N__53182\,
            I => \N__53179\
        );

    \I__12302\ : InMux
    port map (
            O => \N__53179\,
            I => \N__53176\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__53176\,
            I => \N__53172\
        );

    \I__12300\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53169\
        );

    \I__12299\ : Span4Mux_s2_h
    port map (
            O => \N__53172\,
            I => \N__53163\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__53169\,
            I => \N__53163\
        );

    \I__12297\ : InMux
    port map (
            O => \N__53168\,
            I => \N__53160\
        );

    \I__12296\ : Span4Mux_h
    port map (
            O => \N__53163\,
            I => \N__53155\
        );

    \I__12295\ : LocalMux
    port map (
            O => \N__53160\,
            I => \N__53155\
        );

    \I__12294\ : Span4Mux_v
    port map (
            O => \N__53155\,
            I => \N__53152\
        );

    \I__12293\ : Sp12to4
    port map (
            O => \N__53152\,
            I => \N__53149\
        );

    \I__12292\ : Odrv12
    port map (
            O => \N__53149\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__12291\ : InMux
    port map (
            O => \N__53146\,
            I => \N__53143\
        );

    \I__12290\ : LocalMux
    port map (
            O => \N__53143\,
            I => pwm_duty_input_5
        );

    \I__12289\ : InMux
    port map (
            O => \N__53140\,
            I => \N__53137\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__53137\,
            I => \N__53134\
        );

    \I__12287\ : Odrv4
    port map (
            O => \N__53134\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__12286\ : CascadeMux
    port map (
            O => \N__53131\,
            I => \N__53128\
        );

    \I__12285\ : InMux
    port map (
            O => \N__53128\,
            I => \N__53125\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__53125\,
            I => \N__53121\
        );

    \I__12283\ : InMux
    port map (
            O => \N__53124\,
            I => \N__53118\
        );

    \I__12282\ : Odrv4
    port map (
            O => \N__53121\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__12281\ : LocalMux
    port map (
            O => \N__53118\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__12280\ : CascadeMux
    port map (
            O => \N__53113\,
            I => \N__53108\
        );

    \I__12279\ : InMux
    port map (
            O => \N__53112\,
            I => \N__53105\
        );

    \I__12278\ : InMux
    port map (
            O => \N__53111\,
            I => \N__53099\
        );

    \I__12277\ : InMux
    port map (
            O => \N__53108\,
            I => \N__53099\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__53105\,
            I => \N__53096\
        );

    \I__12275\ : InMux
    port map (
            O => \N__53104\,
            I => \N__53093\
        );

    \I__12274\ : LocalMux
    port map (
            O => \N__53099\,
            I => \N__53090\
        );

    \I__12273\ : Span4Mux_v
    port map (
            O => \N__53096\,
            I => \N__53085\
        );

    \I__12272\ : LocalMux
    port map (
            O => \N__53093\,
            I => \N__53085\
        );

    \I__12271\ : Span4Mux_h
    port map (
            O => \N__53090\,
            I => \N__53082\
        );

    \I__12270\ : Span4Mux_h
    port map (
            O => \N__53085\,
            I => \N__53079\
        );

    \I__12269\ : Span4Mux_h
    port map (
            O => \N__53082\,
            I => \N__53076\
        );

    \I__12268\ : Span4Mux_h
    port map (
            O => \N__53079\,
            I => \N__53073\
        );

    \I__12267\ : Span4Mux_h
    port map (
            O => \N__53076\,
            I => \N__53070\
        );

    \I__12266\ : Span4Mux_h
    port map (
            O => \N__53073\,
            I => \N__53067\
        );

    \I__12265\ : Odrv4
    port map (
            O => \N__53070\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__12264\ : Odrv4
    port map (
            O => \N__53067\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__12263\ : InMux
    port map (
            O => \N__53062\,
            I => \N__53059\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__53059\,
            I => pwm_duty_input_4
        );

    \I__12261\ : InMux
    port map (
            O => \N__53056\,
            I => \N__53053\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__53053\,
            I => \N__53048\
        );

    \I__12259\ : InMux
    port map (
            O => \N__53052\,
            I => \N__53045\
        );

    \I__12258\ : InMux
    port map (
            O => \N__53051\,
            I => \N__53042\
        );

    \I__12257\ : Span4Mux_s2_h
    port map (
            O => \N__53048\,
            I => \N__53039\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__53045\,
            I => \N__53034\
        );

    \I__12255\ : LocalMux
    port map (
            O => \N__53042\,
            I => \N__53034\
        );

    \I__12254\ : Span4Mux_v
    port map (
            O => \N__53039\,
            I => \N__53031\
        );

    \I__12253\ : Sp12to4
    port map (
            O => \N__53034\,
            I => \N__53028\
        );

    \I__12252\ : Sp12to4
    port map (
            O => \N__53031\,
            I => \N__53023\
        );

    \I__12251\ : Span12Mux_v
    port map (
            O => \N__53028\,
            I => \N__53023\
        );

    \I__12250\ : Odrv12
    port map (
            O => \N__53023\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__12249\ : InMux
    port map (
            O => \N__53020\,
            I => \N__53017\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__53017\,
            I => pwm_duty_input_7
        );

    \I__12247\ : InMux
    port map (
            O => \N__53014\,
            I => \N__53011\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__53011\,
            I => \N__53008\
        );

    \I__12245\ : Odrv12
    port map (
            O => \N__53008\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__12244\ : InMux
    port map (
            O => \N__53005\,
            I => \N__52998\
        );

    \I__12243\ : InMux
    port map (
            O => \N__53004\,
            I => \N__52998\
        );

    \I__12242\ : InMux
    port map (
            O => \N__53003\,
            I => \N__52995\
        );

    \I__12241\ : LocalMux
    port map (
            O => \N__52998\,
            I => \current_shift_inst.PI_CTRL.N_162\
        );

    \I__12240\ : LocalMux
    port map (
            O => \N__52995\,
            I => \current_shift_inst.PI_CTRL.N_162\
        );

    \I__12239\ : InMux
    port map (
            O => \N__52990\,
            I => \N__52987\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__52987\,
            I => pwm_duty_input_0
        );

    \I__12237\ : InMux
    port map (
            O => \N__52984\,
            I => \N__52980\
        );

    \I__12236\ : InMux
    port map (
            O => \N__52983\,
            I => \N__52977\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__52980\,
            I => \N__52971\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__52977\,
            I => \N__52971\
        );

    \I__12233\ : InMux
    port map (
            O => \N__52976\,
            I => \N__52968\
        );

    \I__12232\ : Span4Mux_v
    port map (
            O => \N__52971\,
            I => \N__52965\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__52968\,
            I => \N__52962\
        );

    \I__12230\ : Span4Mux_h
    port map (
            O => \N__52965\,
            I => \N__52957\
        );

    \I__12229\ : Span4Mux_h
    port map (
            O => \N__52962\,
            I => \N__52957\
        );

    \I__12228\ : Span4Mux_h
    port map (
            O => \N__52957\,
            I => \N__52954\
        );

    \I__12227\ : Span4Mux_h
    port map (
            O => \N__52954\,
            I => \N__52951\
        );

    \I__12226\ : Odrv4
    port map (
            O => \N__52951\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__12225\ : InMux
    port map (
            O => \N__52948\,
            I => \N__52945\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__52945\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__12223\ : InMux
    port map (
            O => \N__52942\,
            I => \N__52939\
        );

    \I__12222\ : LocalMux
    port map (
            O => \N__52939\,
            I => \N__52935\
        );

    \I__12221\ : InMux
    port map (
            O => \N__52938\,
            I => \N__52932\
        );

    \I__12220\ : Odrv4
    port map (
            O => \N__52935\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__12219\ : LocalMux
    port map (
            O => \N__52932\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__12218\ : InMux
    port map (
            O => \N__52927\,
            I => \N__52924\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__52924\,
            I => pwm_duty_input_3
        );

    \I__12216\ : InMux
    port map (
            O => \N__52921\,
            I => \N__52911\
        );

    \I__12215\ : InMux
    port map (
            O => \N__52920\,
            I => \N__52911\
        );

    \I__12214\ : InMux
    port map (
            O => \N__52919\,
            I => \N__52908\
        );

    \I__12213\ : InMux
    port map (
            O => \N__52918\,
            I => \N__52901\
        );

    \I__12212\ : InMux
    port map (
            O => \N__52917\,
            I => \N__52901\
        );

    \I__12211\ : InMux
    port map (
            O => \N__52916\,
            I => \N__52901\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__52911\,
            I => \N__52897\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__52908\,
            I => \N__52894\
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__52901\,
            I => \N__52891\
        );

    \I__12207\ : InMux
    port map (
            O => \N__52900\,
            I => \N__52888\
        );

    \I__12206\ : Span4Mux_v
    port map (
            O => \N__52897\,
            I => \N__52885\
        );

    \I__12205\ : Span4Mux_s3_h
    port map (
            O => \N__52894\,
            I => \N__52882\
        );

    \I__12204\ : Span4Mux_s2_h
    port map (
            O => \N__52891\,
            I => \N__52877\
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__52888\,
            I => \N__52877\
        );

    \I__12202\ : Span4Mux_v
    port map (
            O => \N__52885\,
            I => \N__52871\
        );

    \I__12201\ : Span4Mux_v
    port map (
            O => \N__52882\,
            I => \N__52868\
        );

    \I__12200\ : Span4Mux_v
    port map (
            O => \N__52877\,
            I => \N__52865\
        );

    \I__12199\ : InMux
    port map (
            O => \N__52876\,
            I => \N__52858\
        );

    \I__12198\ : InMux
    port map (
            O => \N__52875\,
            I => \N__52858\
        );

    \I__12197\ : InMux
    port map (
            O => \N__52874\,
            I => \N__52858\
        );

    \I__12196\ : Span4Mux_h
    port map (
            O => \N__52871\,
            I => \N__52855\
        );

    \I__12195\ : Sp12to4
    port map (
            O => \N__52868\,
            I => \N__52852\
        );

    \I__12194\ : Span4Mux_v
    port map (
            O => \N__52865\,
            I => \N__52849\
        );

    \I__12193\ : LocalMux
    port map (
            O => \N__52858\,
            I => \N__52846\
        );

    \I__12192\ : Sp12to4
    port map (
            O => \N__52855\,
            I => \N__52837\
        );

    \I__12191\ : Span12Mux_s7_v
    port map (
            O => \N__52852\,
            I => \N__52837\
        );

    \I__12190\ : Sp12to4
    port map (
            O => \N__52849\,
            I => \N__52837\
        );

    \I__12189\ : Span12Mux_v
    port map (
            O => \N__52846\,
            I => \N__52837\
        );

    \I__12188\ : Odrv12
    port map (
            O => \N__52837\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__12187\ : InMux
    port map (
            O => \N__52834\,
            I => \N__52824\
        );

    \I__12186\ : InMux
    port map (
            O => \N__52833\,
            I => \N__52824\
        );

    \I__12185\ : InMux
    port map (
            O => \N__52832\,
            I => \N__52816\
        );

    \I__12184\ : InMux
    port map (
            O => \N__52831\,
            I => \N__52816\
        );

    \I__12183\ : InMux
    port map (
            O => \N__52830\,
            I => \N__52816\
        );

    \I__12182\ : InMux
    port map (
            O => \N__52829\,
            I => \N__52813\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__52824\,
            I => \N__52810\
        );

    \I__12180\ : InMux
    port map (
            O => \N__52823\,
            I => \N__52807\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__52816\,
            I => \N__52802\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__52813\,
            I => \N__52802\
        );

    \I__12177\ : Span4Mux_s2_h
    port map (
            O => \N__52810\,
            I => \N__52797\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__52807\,
            I => \N__52797\
        );

    \I__12175\ : Span4Mux_v
    port map (
            O => \N__52802\,
            I => \N__52794\
        );

    \I__12174\ : Span4Mux_v
    port map (
            O => \N__52797\,
            I => \N__52791\
        );

    \I__12173\ : Span4Mux_h
    port map (
            O => \N__52794\,
            I => \N__52788\
        );

    \I__12172\ : Span4Mux_h
    port map (
            O => \N__52791\,
            I => \N__52785\
        );

    \I__12171\ : Span4Mux_h
    port map (
            O => \N__52788\,
            I => \N__52782\
        );

    \I__12170\ : Span4Mux_h
    port map (
            O => \N__52785\,
            I => \N__52779\
        );

    \I__12169\ : Odrv4
    port map (
            O => \N__52782\,
            I => \current_shift_inst.PI_CTRL.N_160\
        );

    \I__12168\ : Odrv4
    port map (
            O => \N__52779\,
            I => \current_shift_inst.PI_CTRL.N_160\
        );

    \I__12167\ : CascadeMux
    port map (
            O => \N__52774\,
            I => \N__52771\
        );

    \I__12166\ : InMux
    port map (
            O => \N__52771\,
            I => \N__52767\
        );

    \I__12165\ : InMux
    port map (
            O => \N__52770\,
            I => \N__52764\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__52767\,
            I => \N__52761\
        );

    \I__12163\ : LocalMux
    port map (
            O => \N__52764\,
            I => \N__52758\
        );

    \I__12162\ : Span4Mux_v
    port map (
            O => \N__52761\,
            I => \N__52754\
        );

    \I__12161\ : Span4Mux_h
    port map (
            O => \N__52758\,
            I => \N__52751\
        );

    \I__12160\ : InMux
    port map (
            O => \N__52757\,
            I => \N__52748\
        );

    \I__12159\ : Sp12to4
    port map (
            O => \N__52754\,
            I => \N__52745\
        );

    \I__12158\ : Span4Mux_v
    port map (
            O => \N__52751\,
            I => \N__52742\
        );

    \I__12157\ : LocalMux
    port map (
            O => \N__52748\,
            I => \N__52739\
        );

    \I__12156\ : Span12Mux_s4_h
    port map (
            O => \N__52745\,
            I => \N__52732\
        );

    \I__12155\ : Sp12to4
    port map (
            O => \N__52742\,
            I => \N__52732\
        );

    \I__12154\ : Span12Mux_v
    port map (
            O => \N__52739\,
            I => \N__52732\
        );

    \I__12153\ : Odrv12
    port map (
            O => \N__52732\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__12152\ : CascadeMux
    port map (
            O => \N__52729\,
            I => \N__52723\
        );

    \I__12151\ : CascadeMux
    port map (
            O => \N__52728\,
            I => \N__52719\
        );

    \I__12150\ : InMux
    port map (
            O => \N__52727\,
            I => \N__52715\
        );

    \I__12149\ : InMux
    port map (
            O => \N__52726\,
            I => \N__52710\
        );

    \I__12148\ : InMux
    port map (
            O => \N__52723\,
            I => \N__52710\
        );

    \I__12147\ : InMux
    port map (
            O => \N__52722\,
            I => \N__52705\
        );

    \I__12146\ : InMux
    port map (
            O => \N__52719\,
            I => \N__52705\
        );

    \I__12145\ : CascadeMux
    port map (
            O => \N__52718\,
            I => \N__52702\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__52715\,
            I => \N__52697\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__52710\,
            I => \N__52692\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__52705\,
            I => \N__52692\
        );

    \I__12141\ : InMux
    port map (
            O => \N__52702\,
            I => \N__52687\
        );

    \I__12140\ : InMux
    port map (
            O => \N__52701\,
            I => \N__52687\
        );

    \I__12139\ : InMux
    port map (
            O => \N__52700\,
            I => \N__52684\
        );

    \I__12138\ : Span4Mux_v
    port map (
            O => \N__52697\,
            I => \N__52675\
        );

    \I__12137\ : Span4Mux_v
    port map (
            O => \N__52692\,
            I => \N__52675\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__52687\,
            I => \N__52675\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__52684\,
            I => \N__52675\
        );

    \I__12134\ : Span4Mux_h
    port map (
            O => \N__52675\,
            I => \N__52672\
        );

    \I__12133\ : Span4Mux_v
    port map (
            O => \N__52672\,
            I => \N__52669\
        );

    \I__12132\ : Span4Mux_h
    port map (
            O => \N__52669\,
            I => \N__52666\
        );

    \I__12131\ : Odrv4
    port map (
            O => \N__52666\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\
        );

    \I__12130\ : InMux
    port map (
            O => \N__52663\,
            I => \N__52660\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__52660\,
            I => pwm_duty_input_8
        );

    \I__12128\ : ClkMux
    port map (
            O => \N__52657\,
            I => \N__52297\
        );

    \I__12127\ : ClkMux
    port map (
            O => \N__52656\,
            I => \N__52297\
        );

    \I__12126\ : ClkMux
    port map (
            O => \N__52655\,
            I => \N__52297\
        );

    \I__12125\ : ClkMux
    port map (
            O => \N__52654\,
            I => \N__52297\
        );

    \I__12124\ : ClkMux
    port map (
            O => \N__52653\,
            I => \N__52297\
        );

    \I__12123\ : ClkMux
    port map (
            O => \N__52652\,
            I => \N__52297\
        );

    \I__12122\ : ClkMux
    port map (
            O => \N__52651\,
            I => \N__52297\
        );

    \I__12121\ : ClkMux
    port map (
            O => \N__52650\,
            I => \N__52297\
        );

    \I__12120\ : ClkMux
    port map (
            O => \N__52649\,
            I => \N__52297\
        );

    \I__12119\ : ClkMux
    port map (
            O => \N__52648\,
            I => \N__52297\
        );

    \I__12118\ : ClkMux
    port map (
            O => \N__52647\,
            I => \N__52297\
        );

    \I__12117\ : ClkMux
    port map (
            O => \N__52646\,
            I => \N__52297\
        );

    \I__12116\ : ClkMux
    port map (
            O => \N__52645\,
            I => \N__52297\
        );

    \I__12115\ : ClkMux
    port map (
            O => \N__52644\,
            I => \N__52297\
        );

    \I__12114\ : ClkMux
    port map (
            O => \N__52643\,
            I => \N__52297\
        );

    \I__12113\ : ClkMux
    port map (
            O => \N__52642\,
            I => \N__52297\
        );

    \I__12112\ : ClkMux
    port map (
            O => \N__52641\,
            I => \N__52297\
        );

    \I__12111\ : ClkMux
    port map (
            O => \N__52640\,
            I => \N__52297\
        );

    \I__12110\ : ClkMux
    port map (
            O => \N__52639\,
            I => \N__52297\
        );

    \I__12109\ : ClkMux
    port map (
            O => \N__52638\,
            I => \N__52297\
        );

    \I__12108\ : ClkMux
    port map (
            O => \N__52637\,
            I => \N__52297\
        );

    \I__12107\ : ClkMux
    port map (
            O => \N__52636\,
            I => \N__52297\
        );

    \I__12106\ : ClkMux
    port map (
            O => \N__52635\,
            I => \N__52297\
        );

    \I__12105\ : ClkMux
    port map (
            O => \N__52634\,
            I => \N__52297\
        );

    \I__12104\ : ClkMux
    port map (
            O => \N__52633\,
            I => \N__52297\
        );

    \I__12103\ : ClkMux
    port map (
            O => \N__52632\,
            I => \N__52297\
        );

    \I__12102\ : ClkMux
    port map (
            O => \N__52631\,
            I => \N__52297\
        );

    \I__12101\ : ClkMux
    port map (
            O => \N__52630\,
            I => \N__52297\
        );

    \I__12100\ : ClkMux
    port map (
            O => \N__52629\,
            I => \N__52297\
        );

    \I__12099\ : ClkMux
    port map (
            O => \N__52628\,
            I => \N__52297\
        );

    \I__12098\ : ClkMux
    port map (
            O => \N__52627\,
            I => \N__52297\
        );

    \I__12097\ : ClkMux
    port map (
            O => \N__52626\,
            I => \N__52297\
        );

    \I__12096\ : ClkMux
    port map (
            O => \N__52625\,
            I => \N__52297\
        );

    \I__12095\ : ClkMux
    port map (
            O => \N__52624\,
            I => \N__52297\
        );

    \I__12094\ : ClkMux
    port map (
            O => \N__52623\,
            I => \N__52297\
        );

    \I__12093\ : ClkMux
    port map (
            O => \N__52622\,
            I => \N__52297\
        );

    \I__12092\ : ClkMux
    port map (
            O => \N__52621\,
            I => \N__52297\
        );

    \I__12091\ : ClkMux
    port map (
            O => \N__52620\,
            I => \N__52297\
        );

    \I__12090\ : ClkMux
    port map (
            O => \N__52619\,
            I => \N__52297\
        );

    \I__12089\ : ClkMux
    port map (
            O => \N__52618\,
            I => \N__52297\
        );

    \I__12088\ : ClkMux
    port map (
            O => \N__52617\,
            I => \N__52297\
        );

    \I__12087\ : ClkMux
    port map (
            O => \N__52616\,
            I => \N__52297\
        );

    \I__12086\ : ClkMux
    port map (
            O => \N__52615\,
            I => \N__52297\
        );

    \I__12085\ : ClkMux
    port map (
            O => \N__52614\,
            I => \N__52297\
        );

    \I__12084\ : ClkMux
    port map (
            O => \N__52613\,
            I => \N__52297\
        );

    \I__12083\ : ClkMux
    port map (
            O => \N__52612\,
            I => \N__52297\
        );

    \I__12082\ : ClkMux
    port map (
            O => \N__52611\,
            I => \N__52297\
        );

    \I__12081\ : ClkMux
    port map (
            O => \N__52610\,
            I => \N__52297\
        );

    \I__12080\ : ClkMux
    port map (
            O => \N__52609\,
            I => \N__52297\
        );

    \I__12079\ : ClkMux
    port map (
            O => \N__52608\,
            I => \N__52297\
        );

    \I__12078\ : ClkMux
    port map (
            O => \N__52607\,
            I => \N__52297\
        );

    \I__12077\ : ClkMux
    port map (
            O => \N__52606\,
            I => \N__52297\
        );

    \I__12076\ : ClkMux
    port map (
            O => \N__52605\,
            I => \N__52297\
        );

    \I__12075\ : ClkMux
    port map (
            O => \N__52604\,
            I => \N__52297\
        );

    \I__12074\ : ClkMux
    port map (
            O => \N__52603\,
            I => \N__52297\
        );

    \I__12073\ : ClkMux
    port map (
            O => \N__52602\,
            I => \N__52297\
        );

    \I__12072\ : ClkMux
    port map (
            O => \N__52601\,
            I => \N__52297\
        );

    \I__12071\ : ClkMux
    port map (
            O => \N__52600\,
            I => \N__52297\
        );

    \I__12070\ : ClkMux
    port map (
            O => \N__52599\,
            I => \N__52297\
        );

    \I__12069\ : ClkMux
    port map (
            O => \N__52598\,
            I => \N__52297\
        );

    \I__12068\ : ClkMux
    port map (
            O => \N__52597\,
            I => \N__52297\
        );

    \I__12067\ : ClkMux
    port map (
            O => \N__52596\,
            I => \N__52297\
        );

    \I__12066\ : ClkMux
    port map (
            O => \N__52595\,
            I => \N__52297\
        );

    \I__12065\ : ClkMux
    port map (
            O => \N__52594\,
            I => \N__52297\
        );

    \I__12064\ : ClkMux
    port map (
            O => \N__52593\,
            I => \N__52297\
        );

    \I__12063\ : ClkMux
    port map (
            O => \N__52592\,
            I => \N__52297\
        );

    \I__12062\ : ClkMux
    port map (
            O => \N__52591\,
            I => \N__52297\
        );

    \I__12061\ : ClkMux
    port map (
            O => \N__52590\,
            I => \N__52297\
        );

    \I__12060\ : ClkMux
    port map (
            O => \N__52589\,
            I => \N__52297\
        );

    \I__12059\ : ClkMux
    port map (
            O => \N__52588\,
            I => \N__52297\
        );

    \I__12058\ : ClkMux
    port map (
            O => \N__52587\,
            I => \N__52297\
        );

    \I__12057\ : ClkMux
    port map (
            O => \N__52586\,
            I => \N__52297\
        );

    \I__12056\ : ClkMux
    port map (
            O => \N__52585\,
            I => \N__52297\
        );

    \I__12055\ : ClkMux
    port map (
            O => \N__52584\,
            I => \N__52297\
        );

    \I__12054\ : ClkMux
    port map (
            O => \N__52583\,
            I => \N__52297\
        );

    \I__12053\ : ClkMux
    port map (
            O => \N__52582\,
            I => \N__52297\
        );

    \I__12052\ : ClkMux
    port map (
            O => \N__52581\,
            I => \N__52297\
        );

    \I__12051\ : ClkMux
    port map (
            O => \N__52580\,
            I => \N__52297\
        );

    \I__12050\ : ClkMux
    port map (
            O => \N__52579\,
            I => \N__52297\
        );

    \I__12049\ : ClkMux
    port map (
            O => \N__52578\,
            I => \N__52297\
        );

    \I__12048\ : ClkMux
    port map (
            O => \N__52577\,
            I => \N__52297\
        );

    \I__12047\ : ClkMux
    port map (
            O => \N__52576\,
            I => \N__52297\
        );

    \I__12046\ : ClkMux
    port map (
            O => \N__52575\,
            I => \N__52297\
        );

    \I__12045\ : ClkMux
    port map (
            O => \N__52574\,
            I => \N__52297\
        );

    \I__12044\ : ClkMux
    port map (
            O => \N__52573\,
            I => \N__52297\
        );

    \I__12043\ : ClkMux
    port map (
            O => \N__52572\,
            I => \N__52297\
        );

    \I__12042\ : ClkMux
    port map (
            O => \N__52571\,
            I => \N__52297\
        );

    \I__12041\ : ClkMux
    port map (
            O => \N__52570\,
            I => \N__52297\
        );

    \I__12040\ : ClkMux
    port map (
            O => \N__52569\,
            I => \N__52297\
        );

    \I__12039\ : ClkMux
    port map (
            O => \N__52568\,
            I => \N__52297\
        );

    \I__12038\ : ClkMux
    port map (
            O => \N__52567\,
            I => \N__52297\
        );

    \I__12037\ : ClkMux
    port map (
            O => \N__52566\,
            I => \N__52297\
        );

    \I__12036\ : ClkMux
    port map (
            O => \N__52565\,
            I => \N__52297\
        );

    \I__12035\ : ClkMux
    port map (
            O => \N__52564\,
            I => \N__52297\
        );

    \I__12034\ : ClkMux
    port map (
            O => \N__52563\,
            I => \N__52297\
        );

    \I__12033\ : ClkMux
    port map (
            O => \N__52562\,
            I => \N__52297\
        );

    \I__12032\ : ClkMux
    port map (
            O => \N__52561\,
            I => \N__52297\
        );

    \I__12031\ : ClkMux
    port map (
            O => \N__52560\,
            I => \N__52297\
        );

    \I__12030\ : ClkMux
    port map (
            O => \N__52559\,
            I => \N__52297\
        );

    \I__12029\ : ClkMux
    port map (
            O => \N__52558\,
            I => \N__52297\
        );

    \I__12028\ : ClkMux
    port map (
            O => \N__52557\,
            I => \N__52297\
        );

    \I__12027\ : ClkMux
    port map (
            O => \N__52556\,
            I => \N__52297\
        );

    \I__12026\ : ClkMux
    port map (
            O => \N__52555\,
            I => \N__52297\
        );

    \I__12025\ : ClkMux
    port map (
            O => \N__52554\,
            I => \N__52297\
        );

    \I__12024\ : ClkMux
    port map (
            O => \N__52553\,
            I => \N__52297\
        );

    \I__12023\ : ClkMux
    port map (
            O => \N__52552\,
            I => \N__52297\
        );

    \I__12022\ : ClkMux
    port map (
            O => \N__52551\,
            I => \N__52297\
        );

    \I__12021\ : ClkMux
    port map (
            O => \N__52550\,
            I => \N__52297\
        );

    \I__12020\ : ClkMux
    port map (
            O => \N__52549\,
            I => \N__52297\
        );

    \I__12019\ : ClkMux
    port map (
            O => \N__52548\,
            I => \N__52297\
        );

    \I__12018\ : ClkMux
    port map (
            O => \N__52547\,
            I => \N__52297\
        );

    \I__12017\ : ClkMux
    port map (
            O => \N__52546\,
            I => \N__52297\
        );

    \I__12016\ : ClkMux
    port map (
            O => \N__52545\,
            I => \N__52297\
        );

    \I__12015\ : ClkMux
    port map (
            O => \N__52544\,
            I => \N__52297\
        );

    \I__12014\ : ClkMux
    port map (
            O => \N__52543\,
            I => \N__52297\
        );

    \I__12013\ : ClkMux
    port map (
            O => \N__52542\,
            I => \N__52297\
        );

    \I__12012\ : ClkMux
    port map (
            O => \N__52541\,
            I => \N__52297\
        );

    \I__12011\ : ClkMux
    port map (
            O => \N__52540\,
            I => \N__52297\
        );

    \I__12010\ : ClkMux
    port map (
            O => \N__52539\,
            I => \N__52297\
        );

    \I__12009\ : ClkMux
    port map (
            O => \N__52538\,
            I => \N__52297\
        );

    \I__12008\ : GlobalMux
    port map (
            O => \N__52297\,
            I => clk_100mhz_0
        );

    \I__12007\ : InMux
    port map (
            O => \N__52294\,
            I => \N__52287\
        );

    \I__12006\ : InMux
    port map (
            O => \N__52293\,
            I => \N__52284\
        );

    \I__12005\ : InMux
    port map (
            O => \N__52292\,
            I => \N__52281\
        );

    \I__12004\ : InMux
    port map (
            O => \N__52291\,
            I => \N__52278\
        );

    \I__12003\ : InMux
    port map (
            O => \N__52290\,
            I => \N__52275\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__52287\,
            I => \N__52272\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__52284\,
            I => \N__52226\
        );

    \I__12000\ : LocalMux
    port map (
            O => \N__52281\,
            I => \N__52203\
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__52278\,
            I => \N__52200\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__52275\,
            I => \N__52184\
        );

    \I__11997\ : Glb2LocalMux
    port map (
            O => \N__52272\,
            I => \N__51973\
        );

    \I__11996\ : SRMux
    port map (
            O => \N__52271\,
            I => \N__51973\
        );

    \I__11995\ : SRMux
    port map (
            O => \N__52270\,
            I => \N__51973\
        );

    \I__11994\ : SRMux
    port map (
            O => \N__52269\,
            I => \N__51973\
        );

    \I__11993\ : SRMux
    port map (
            O => \N__52268\,
            I => \N__51973\
        );

    \I__11992\ : SRMux
    port map (
            O => \N__52267\,
            I => \N__51973\
        );

    \I__11991\ : SRMux
    port map (
            O => \N__52266\,
            I => \N__51973\
        );

    \I__11990\ : SRMux
    port map (
            O => \N__52265\,
            I => \N__51973\
        );

    \I__11989\ : SRMux
    port map (
            O => \N__52264\,
            I => \N__51973\
        );

    \I__11988\ : SRMux
    port map (
            O => \N__52263\,
            I => \N__51973\
        );

    \I__11987\ : SRMux
    port map (
            O => \N__52262\,
            I => \N__51973\
        );

    \I__11986\ : SRMux
    port map (
            O => \N__52261\,
            I => \N__51973\
        );

    \I__11985\ : SRMux
    port map (
            O => \N__52260\,
            I => \N__51973\
        );

    \I__11984\ : SRMux
    port map (
            O => \N__52259\,
            I => \N__51973\
        );

    \I__11983\ : SRMux
    port map (
            O => \N__52258\,
            I => \N__51973\
        );

    \I__11982\ : SRMux
    port map (
            O => \N__52257\,
            I => \N__51973\
        );

    \I__11981\ : SRMux
    port map (
            O => \N__52256\,
            I => \N__51973\
        );

    \I__11980\ : SRMux
    port map (
            O => \N__52255\,
            I => \N__51973\
        );

    \I__11979\ : SRMux
    port map (
            O => \N__52254\,
            I => \N__51973\
        );

    \I__11978\ : SRMux
    port map (
            O => \N__52253\,
            I => \N__51973\
        );

    \I__11977\ : SRMux
    port map (
            O => \N__52252\,
            I => \N__51973\
        );

    \I__11976\ : SRMux
    port map (
            O => \N__52251\,
            I => \N__51973\
        );

    \I__11975\ : SRMux
    port map (
            O => \N__52250\,
            I => \N__51973\
        );

    \I__11974\ : SRMux
    port map (
            O => \N__52249\,
            I => \N__51973\
        );

    \I__11973\ : SRMux
    port map (
            O => \N__52248\,
            I => \N__51973\
        );

    \I__11972\ : SRMux
    port map (
            O => \N__52247\,
            I => \N__51973\
        );

    \I__11971\ : SRMux
    port map (
            O => \N__52246\,
            I => \N__51973\
        );

    \I__11970\ : SRMux
    port map (
            O => \N__52245\,
            I => \N__51973\
        );

    \I__11969\ : SRMux
    port map (
            O => \N__52244\,
            I => \N__51973\
        );

    \I__11968\ : SRMux
    port map (
            O => \N__52243\,
            I => \N__51973\
        );

    \I__11967\ : SRMux
    port map (
            O => \N__52242\,
            I => \N__51973\
        );

    \I__11966\ : SRMux
    port map (
            O => \N__52241\,
            I => \N__51973\
        );

    \I__11965\ : SRMux
    port map (
            O => \N__52240\,
            I => \N__51973\
        );

    \I__11964\ : SRMux
    port map (
            O => \N__52239\,
            I => \N__51973\
        );

    \I__11963\ : SRMux
    port map (
            O => \N__52238\,
            I => \N__51973\
        );

    \I__11962\ : SRMux
    port map (
            O => \N__52237\,
            I => \N__51973\
        );

    \I__11961\ : SRMux
    port map (
            O => \N__52236\,
            I => \N__51973\
        );

    \I__11960\ : SRMux
    port map (
            O => \N__52235\,
            I => \N__51973\
        );

    \I__11959\ : SRMux
    port map (
            O => \N__52234\,
            I => \N__51973\
        );

    \I__11958\ : SRMux
    port map (
            O => \N__52233\,
            I => \N__51973\
        );

    \I__11957\ : SRMux
    port map (
            O => \N__52232\,
            I => \N__51973\
        );

    \I__11956\ : SRMux
    port map (
            O => \N__52231\,
            I => \N__51973\
        );

    \I__11955\ : SRMux
    port map (
            O => \N__52230\,
            I => \N__51973\
        );

    \I__11954\ : SRMux
    port map (
            O => \N__52229\,
            I => \N__51973\
        );

    \I__11953\ : Glb2LocalMux
    port map (
            O => \N__52226\,
            I => \N__51973\
        );

    \I__11952\ : SRMux
    port map (
            O => \N__52225\,
            I => \N__51973\
        );

    \I__11951\ : SRMux
    port map (
            O => \N__52224\,
            I => \N__51973\
        );

    \I__11950\ : SRMux
    port map (
            O => \N__52223\,
            I => \N__51973\
        );

    \I__11949\ : SRMux
    port map (
            O => \N__52222\,
            I => \N__51973\
        );

    \I__11948\ : SRMux
    port map (
            O => \N__52221\,
            I => \N__51973\
        );

    \I__11947\ : SRMux
    port map (
            O => \N__52220\,
            I => \N__51973\
        );

    \I__11946\ : SRMux
    port map (
            O => \N__52219\,
            I => \N__51973\
        );

    \I__11945\ : SRMux
    port map (
            O => \N__52218\,
            I => \N__51973\
        );

    \I__11944\ : SRMux
    port map (
            O => \N__52217\,
            I => \N__51973\
        );

    \I__11943\ : SRMux
    port map (
            O => \N__52216\,
            I => \N__51973\
        );

    \I__11942\ : SRMux
    port map (
            O => \N__52215\,
            I => \N__51973\
        );

    \I__11941\ : SRMux
    port map (
            O => \N__52214\,
            I => \N__51973\
        );

    \I__11940\ : SRMux
    port map (
            O => \N__52213\,
            I => \N__51973\
        );

    \I__11939\ : SRMux
    port map (
            O => \N__52212\,
            I => \N__51973\
        );

    \I__11938\ : SRMux
    port map (
            O => \N__52211\,
            I => \N__51973\
        );

    \I__11937\ : SRMux
    port map (
            O => \N__52210\,
            I => \N__51973\
        );

    \I__11936\ : SRMux
    port map (
            O => \N__52209\,
            I => \N__51973\
        );

    \I__11935\ : SRMux
    port map (
            O => \N__52208\,
            I => \N__51973\
        );

    \I__11934\ : SRMux
    port map (
            O => \N__52207\,
            I => \N__51973\
        );

    \I__11933\ : SRMux
    port map (
            O => \N__52206\,
            I => \N__51973\
        );

    \I__11932\ : Glb2LocalMux
    port map (
            O => \N__52203\,
            I => \N__51973\
        );

    \I__11931\ : Glb2LocalMux
    port map (
            O => \N__52200\,
            I => \N__51973\
        );

    \I__11930\ : SRMux
    port map (
            O => \N__52199\,
            I => \N__51973\
        );

    \I__11929\ : SRMux
    port map (
            O => \N__52198\,
            I => \N__51973\
        );

    \I__11928\ : SRMux
    port map (
            O => \N__52197\,
            I => \N__51973\
        );

    \I__11927\ : SRMux
    port map (
            O => \N__52196\,
            I => \N__51973\
        );

    \I__11926\ : SRMux
    port map (
            O => \N__52195\,
            I => \N__51973\
        );

    \I__11925\ : SRMux
    port map (
            O => \N__52194\,
            I => \N__51973\
        );

    \I__11924\ : SRMux
    port map (
            O => \N__52193\,
            I => \N__51973\
        );

    \I__11923\ : SRMux
    port map (
            O => \N__52192\,
            I => \N__51973\
        );

    \I__11922\ : SRMux
    port map (
            O => \N__52191\,
            I => \N__51973\
        );

    \I__11921\ : SRMux
    port map (
            O => \N__52190\,
            I => \N__51973\
        );

    \I__11920\ : SRMux
    port map (
            O => \N__52189\,
            I => \N__51973\
        );

    \I__11919\ : SRMux
    port map (
            O => \N__52188\,
            I => \N__51973\
        );

    \I__11918\ : SRMux
    port map (
            O => \N__52187\,
            I => \N__51973\
        );

    \I__11917\ : Glb2LocalMux
    port map (
            O => \N__52184\,
            I => \N__51973\
        );

    \I__11916\ : SRMux
    port map (
            O => \N__52183\,
            I => \N__51973\
        );

    \I__11915\ : SRMux
    port map (
            O => \N__52182\,
            I => \N__51973\
        );

    \I__11914\ : SRMux
    port map (
            O => \N__52181\,
            I => \N__51973\
        );

    \I__11913\ : SRMux
    port map (
            O => \N__52180\,
            I => \N__51973\
        );

    \I__11912\ : SRMux
    port map (
            O => \N__52179\,
            I => \N__51973\
        );

    \I__11911\ : SRMux
    port map (
            O => \N__52178\,
            I => \N__51973\
        );

    \I__11910\ : SRMux
    port map (
            O => \N__52177\,
            I => \N__51973\
        );

    \I__11909\ : SRMux
    port map (
            O => \N__52176\,
            I => \N__51973\
        );

    \I__11908\ : SRMux
    port map (
            O => \N__52175\,
            I => \N__51973\
        );

    \I__11907\ : SRMux
    port map (
            O => \N__52174\,
            I => \N__51973\
        );

    \I__11906\ : SRMux
    port map (
            O => \N__52173\,
            I => \N__51973\
        );

    \I__11905\ : SRMux
    port map (
            O => \N__52172\,
            I => \N__51973\
        );

    \I__11904\ : SRMux
    port map (
            O => \N__52171\,
            I => \N__51973\
        );

    \I__11903\ : SRMux
    port map (
            O => \N__52170\,
            I => \N__51973\
        );

    \I__11902\ : SRMux
    port map (
            O => \N__52169\,
            I => \N__51973\
        );

    \I__11901\ : SRMux
    port map (
            O => \N__52168\,
            I => \N__51973\
        );

    \I__11900\ : GlobalMux
    port map (
            O => \N__51973\,
            I => \N__51970\
        );

    \I__11899\ : gio2CtrlBuf
    port map (
            O => \N__51970\,
            I => reset_c_g
        );

    \I__11898\ : InMux
    port map (
            O => \N__51967\,
            I => \N__51964\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__51964\,
            I => \current_shift_inst.PI_CTRL.N_145\
        );

    \I__11896\ : CascadeMux
    port map (
            O => \N__51961\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__11895\ : CascadeMux
    port map (
            O => \N__51958\,
            I => \N__51955\
        );

    \I__11894\ : InMux
    port map (
            O => \N__51955\,
            I => \N__51952\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__51952\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__11892\ : InMux
    port map (
            O => \N__51949\,
            I => \N__51946\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__51946\,
            I => \N__51942\
        );

    \I__11890\ : InMux
    port map (
            O => \N__51945\,
            I => \N__51939\
        );

    \I__11889\ : Span12Mux_s8_v
    port map (
            O => \N__51942\,
            I => \N__51936\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__51939\,
            I => \N__51933\
        );

    \I__11887\ : Span12Mux_h
    port map (
            O => \N__51936\,
            I => \N__51930\
        );

    \I__11886\ : Sp12to4
    port map (
            O => \N__51933\,
            I => \N__51925\
        );

    \I__11885\ : Span12Mux_h
    port map (
            O => \N__51930\,
            I => \N__51925\
        );

    \I__11884\ : Odrv12
    port map (
            O => \N__51925\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__11883\ : InMux
    port map (
            O => \N__51922\,
            I => \N__51919\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__51919\,
            I => \N__51916\
        );

    \I__11881\ : Span12Mux_v
    port map (
            O => \N__51916\,
            I => \N__51913\
        );

    \I__11880\ : Span12Mux_h
    port map (
            O => \N__51913\,
            I => \N__51910\
        );

    \I__11879\ : Span12Mux_h
    port map (
            O => \N__51910\,
            I => \N__51907\
        );

    \I__11878\ : Odrv12
    port map (
            O => \N__51907\,
            I => \pwm_generator_inst.un3_threshold_iZ0\
        );

    \I__11877\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51900\
        );

    \I__11876\ : InMux
    port map (
            O => \N__51903\,
            I => \N__51897\
        );

    \I__11875\ : LocalMux
    port map (
            O => \N__51900\,
            I => \N__51894\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__51897\,
            I => \N__51891\
        );

    \I__11873\ : Span4Mux_v
    port map (
            O => \N__51894\,
            I => \N__51887\
        );

    \I__11872\ : Span4Mux_v
    port map (
            O => \N__51891\,
            I => \N__51884\
        );

    \I__11871\ : InMux
    port map (
            O => \N__51890\,
            I => \N__51881\
        );

    \I__11870\ : Sp12to4
    port map (
            O => \N__51887\,
            I => \N__51874\
        );

    \I__11869\ : Sp12to4
    port map (
            O => \N__51884\,
            I => \N__51874\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__51881\,
            I => \N__51874\
        );

    \I__11867\ : Span12Mux_h
    port map (
            O => \N__51874\,
            I => \N__51871\
        );

    \I__11866\ : Odrv12
    port map (
            O => \N__51871\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__11865\ : InMux
    port map (
            O => \N__51868\,
            I => \N__51865\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__51865\,
            I => \N__51862\
        );

    \I__11863\ : Odrv4
    port map (
            O => \N__51862\,
            I => pwm_duty_input_9
        );

    \I__11862\ : InMux
    port map (
            O => \N__51859\,
            I => \N__51827\
        );

    \I__11861\ : InMux
    port map (
            O => \N__51858\,
            I => \N__51827\
        );

    \I__11860\ : InMux
    port map (
            O => \N__51857\,
            I => \N__51827\
        );

    \I__11859\ : InMux
    port map (
            O => \N__51856\,
            I => \N__51827\
        );

    \I__11858\ : InMux
    port map (
            O => \N__51855\,
            I => \N__51827\
        );

    \I__11857\ : InMux
    port map (
            O => \N__51854\,
            I => \N__51827\
        );

    \I__11856\ : InMux
    port map (
            O => \N__51853\,
            I => \N__51827\
        );

    \I__11855\ : InMux
    port map (
            O => \N__51852\,
            I => \N__51827\
        );

    \I__11854\ : InMux
    port map (
            O => \N__51851\,
            I => \N__51810\
        );

    \I__11853\ : InMux
    port map (
            O => \N__51850\,
            I => \N__51810\
        );

    \I__11852\ : InMux
    port map (
            O => \N__51849\,
            I => \N__51810\
        );

    \I__11851\ : InMux
    port map (
            O => \N__51848\,
            I => \N__51810\
        );

    \I__11850\ : InMux
    port map (
            O => \N__51847\,
            I => \N__51810\
        );

    \I__11849\ : InMux
    port map (
            O => \N__51846\,
            I => \N__51810\
        );

    \I__11848\ : InMux
    port map (
            O => \N__51845\,
            I => \N__51810\
        );

    \I__11847\ : InMux
    port map (
            O => \N__51844\,
            I => \N__51810\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__51827\,
            I => \N__51805\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__51810\,
            I => \N__51805\
        );

    \I__11844\ : Span12Mux_v
    port map (
            O => \N__51805\,
            I => \N__51802\
        );

    \I__11843\ : Span12Mux_h
    port map (
            O => \N__51802\,
            I => \N__51794\
        );

    \I__11842\ : InMux
    port map (
            O => \N__51801\,
            I => \N__51789\
        );

    \I__11841\ : InMux
    port map (
            O => \N__51800\,
            I => \N__51789\
        );

    \I__11840\ : InMux
    port map (
            O => \N__51799\,
            I => \N__51782\
        );

    \I__11839\ : InMux
    port map (
            O => \N__51798\,
            I => \N__51782\
        );

    \I__11838\ : InMux
    port map (
            O => \N__51797\,
            I => \N__51782\
        );

    \I__11837\ : Span12Mux_h
    port map (
            O => \N__51794\,
            I => \N__51779\
        );

    \I__11836\ : LocalMux
    port map (
            O => \N__51789\,
            I => \N__51774\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__51782\,
            I => \N__51774\
        );

    \I__11834\ : Odrv12
    port map (
            O => \N__51779\,
            I => pwm_duty_input_10
        );

    \I__11833\ : Odrv4
    port map (
            O => \N__51774\,
            I => pwm_duty_input_10
        );

    \I__11832\ : InMux
    port map (
            O => \N__51769\,
            I => \N__51766\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__51766\,
            I => \N__51763\
        );

    \I__11830\ : Span4Mux_h
    port map (
            O => \N__51763\,
            I => \N__51760\
        );

    \I__11829\ : Span4Mux_v
    port map (
            O => \N__51760\,
            I => \N__51757\
        );

    \I__11828\ : Sp12to4
    port map (
            O => \N__51757\,
            I => \N__51754\
        );

    \I__11827\ : Odrv12
    port map (
            O => \N__51754\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__11826\ : InMux
    port map (
            O => \N__51751\,
            I => \N__51748\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__51748\,
            I => \N__51745\
        );

    \I__11824\ : Odrv4
    port map (
            O => \N__51745\,
            I => pwm_duty_input_1
        );

    \I__11823\ : InMux
    port map (
            O => \N__51742\,
            I => \N__51739\
        );

    \I__11822\ : LocalMux
    port map (
            O => \N__51739\,
            I => \N__51736\
        );

    \I__11821\ : Span12Mux_v
    port map (
            O => \N__51736\,
            I => \N__51733\
        );

    \I__11820\ : Span12Mux_h
    port map (
            O => \N__51733\,
            I => \N__51730\
        );

    \I__11819\ : Odrv12
    port map (
            O => \N__51730\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__11818\ : InMux
    port map (
            O => \N__51727\,
            I => \N__51724\
        );

    \I__11817\ : LocalMux
    port map (
            O => \N__51724\,
            I => \N__51721\
        );

    \I__11816\ : Span4Mux_v
    port map (
            O => \N__51721\,
            I => \N__51718\
        );

    \I__11815\ : Odrv4
    port map (
            O => \N__51718\,
            I => pwm_duty_input_2
        );

    \I__11814\ : CascadeMux
    port map (
            O => \N__51715\,
            I => \N__51712\
        );

    \I__11813\ : InMux
    port map (
            O => \N__51712\,
            I => \N__51708\
        );

    \I__11812\ : CascadeMux
    port map (
            O => \N__51711\,
            I => \N__51705\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__51708\,
            I => \N__51701\
        );

    \I__11810\ : InMux
    port map (
            O => \N__51705\,
            I => \N__51698\
        );

    \I__11809\ : InMux
    port map (
            O => \N__51704\,
            I => \N__51695\
        );

    \I__11808\ : Span4Mux_v
    port map (
            O => \N__51701\,
            I => \N__51688\
        );

    \I__11807\ : LocalMux
    port map (
            O => \N__51698\,
            I => \N__51688\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__51695\,
            I => \N__51688\
        );

    \I__11805\ : Span4Mux_h
    port map (
            O => \N__51688\,
            I => \N__51685\
        );

    \I__11804\ : Span4Mux_h
    port map (
            O => \N__51685\,
            I => \N__51682\
        );

    \I__11803\ : Span4Mux_h
    port map (
            O => \N__51682\,
            I => \N__51679\
        );

    \I__11802\ : Odrv4
    port map (
            O => \N__51679\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__11801\ : InMux
    port map (
            O => \N__51676\,
            I => \N__51673\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__51673\,
            I => \N__51670\
        );

    \I__11799\ : Odrv4
    port map (
            O => \N__51670\,
            I => pwm_duty_input_6
        );

    \I__11798\ : InMux
    port map (
            O => \N__51667\,
            I => \N__51664\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__51664\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__11796\ : CascadeMux
    port map (
            O => \N__51661\,
            I => \N__51656\
        );

    \I__11795\ : CascadeMux
    port map (
            O => \N__51660\,
            I => \N__51653\
        );

    \I__11794\ : CascadeMux
    port map (
            O => \N__51659\,
            I => \N__51650\
        );

    \I__11793\ : InMux
    port map (
            O => \N__51656\,
            I => \N__51635\
        );

    \I__11792\ : InMux
    port map (
            O => \N__51653\,
            I => \N__51635\
        );

    \I__11791\ : InMux
    port map (
            O => \N__51650\,
            I => \N__51635\
        );

    \I__11790\ : CascadeMux
    port map (
            O => \N__51649\,
            I => \N__51632\
        );

    \I__11789\ : CascadeMux
    port map (
            O => \N__51648\,
            I => \N__51629\
        );

    \I__11788\ : CascadeMux
    port map (
            O => \N__51647\,
            I => \N__51626\
        );

    \I__11787\ : CascadeMux
    port map (
            O => \N__51646\,
            I => \N__51623\
        );

    \I__11786\ : InMux
    port map (
            O => \N__51645\,
            I => \N__51616\
        );

    \I__11785\ : InMux
    port map (
            O => \N__51644\,
            I => \N__51611\
        );

    \I__11784\ : InMux
    port map (
            O => \N__51643\,
            I => \N__51611\
        );

    \I__11783\ : InMux
    port map (
            O => \N__51642\,
            I => \N__51608\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__51635\,
            I => \N__51601\
        );

    \I__11781\ : InMux
    port map (
            O => \N__51632\,
            I => \N__51592\
        );

    \I__11780\ : InMux
    port map (
            O => \N__51629\,
            I => \N__51592\
        );

    \I__11779\ : InMux
    port map (
            O => \N__51626\,
            I => \N__51592\
        );

    \I__11778\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51592\
        );

    \I__11777\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51574\
        );

    \I__11776\ : InMux
    port map (
            O => \N__51621\,
            I => \N__51569\
        );

    \I__11775\ : InMux
    port map (
            O => \N__51620\,
            I => \N__51569\
        );

    \I__11774\ : InMux
    port map (
            O => \N__51619\,
            I => \N__51566\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__51616\,
            I => \N__51559\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__51611\,
            I => \N__51559\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__51608\,
            I => \N__51559\
        );

    \I__11770\ : CascadeMux
    port map (
            O => \N__51607\,
            I => \N__51556\
        );

    \I__11769\ : CascadeMux
    port map (
            O => \N__51606\,
            I => \N__51553\
        );

    \I__11768\ : CascadeMux
    port map (
            O => \N__51605\,
            I => \N__51550\
        );

    \I__11767\ : CascadeMux
    port map (
            O => \N__51604\,
            I => \N__51547\
        );

    \I__11766\ : Span4Mux_v
    port map (
            O => \N__51601\,
            I => \N__51544\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__51592\,
            I => \N__51541\
        );

    \I__11764\ : CascadeMux
    port map (
            O => \N__51591\,
            I => \N__51538\
        );

    \I__11763\ : CascadeMux
    port map (
            O => \N__51590\,
            I => \N__51535\
        );

    \I__11762\ : CascadeMux
    port map (
            O => \N__51589\,
            I => \N__51532\
        );

    \I__11761\ : CascadeMux
    port map (
            O => \N__51588\,
            I => \N__51529\
        );

    \I__11760\ : CascadeMux
    port map (
            O => \N__51587\,
            I => \N__51526\
        );

    \I__11759\ : CascadeMux
    port map (
            O => \N__51586\,
            I => \N__51523\
        );

    \I__11758\ : CascadeMux
    port map (
            O => \N__51585\,
            I => \N__51520\
        );

    \I__11757\ : CascadeMux
    port map (
            O => \N__51584\,
            I => \N__51517\
        );

    \I__11756\ : CascadeMux
    port map (
            O => \N__51583\,
            I => \N__51514\
        );

    \I__11755\ : CascadeMux
    port map (
            O => \N__51582\,
            I => \N__51511\
        );

    \I__11754\ : CascadeMux
    port map (
            O => \N__51581\,
            I => \N__51508\
        );

    \I__11753\ : CascadeMux
    port map (
            O => \N__51580\,
            I => \N__51505\
        );

    \I__11752\ : InMux
    port map (
            O => \N__51579\,
            I => \N__51489\
        );

    \I__11751\ : InMux
    port map (
            O => \N__51578\,
            I => \N__51489\
        );

    \I__11750\ : InMux
    port map (
            O => \N__51577\,
            I => \N__51486\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__51574\,
            I => \N__51479\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__51569\,
            I => \N__51479\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51566\,
            I => \N__51479\
        );

    \I__11746\ : Span4Mux_v
    port map (
            O => \N__51559\,
            I => \N__51476\
        );

    \I__11745\ : InMux
    port map (
            O => \N__51556\,
            I => \N__51454\
        );

    \I__11744\ : InMux
    port map (
            O => \N__51553\,
            I => \N__51454\
        );

    \I__11743\ : InMux
    port map (
            O => \N__51550\,
            I => \N__51454\
        );

    \I__11742\ : InMux
    port map (
            O => \N__51547\,
            I => \N__51454\
        );

    \I__11741\ : Span4Mux_h
    port map (
            O => \N__51544\,
            I => \N__51449\
        );

    \I__11740\ : Span4Mux_v
    port map (
            O => \N__51541\,
            I => \N__51449\
        );

    \I__11739\ : InMux
    port map (
            O => \N__51538\,
            I => \N__51440\
        );

    \I__11738\ : InMux
    port map (
            O => \N__51535\,
            I => \N__51440\
        );

    \I__11737\ : InMux
    port map (
            O => \N__51532\,
            I => \N__51440\
        );

    \I__11736\ : InMux
    port map (
            O => \N__51529\,
            I => \N__51440\
        );

    \I__11735\ : InMux
    port map (
            O => \N__51526\,
            I => \N__51431\
        );

    \I__11734\ : InMux
    port map (
            O => \N__51523\,
            I => \N__51431\
        );

    \I__11733\ : InMux
    port map (
            O => \N__51520\,
            I => \N__51431\
        );

    \I__11732\ : InMux
    port map (
            O => \N__51517\,
            I => \N__51431\
        );

    \I__11731\ : InMux
    port map (
            O => \N__51514\,
            I => \N__51422\
        );

    \I__11730\ : InMux
    port map (
            O => \N__51511\,
            I => \N__51422\
        );

    \I__11729\ : InMux
    port map (
            O => \N__51508\,
            I => \N__51422\
        );

    \I__11728\ : InMux
    port map (
            O => \N__51505\,
            I => \N__51422\
        );

    \I__11727\ : CascadeMux
    port map (
            O => \N__51504\,
            I => \N__51414\
        );

    \I__11726\ : CascadeMux
    port map (
            O => \N__51503\,
            I => \N__51410\
        );

    \I__11725\ : CascadeMux
    port map (
            O => \N__51502\,
            I => \N__51406\
        );

    \I__11724\ : CascadeMux
    port map (
            O => \N__51501\,
            I => \N__51402\
        );

    \I__11723\ : CascadeMux
    port map (
            O => \N__51500\,
            I => \N__51398\
        );

    \I__11722\ : CascadeMux
    port map (
            O => \N__51499\,
            I => \N__51394\
        );

    \I__11721\ : CascadeMux
    port map (
            O => \N__51498\,
            I => \N__51390\
        );

    \I__11720\ : CascadeMux
    port map (
            O => \N__51497\,
            I => \N__51383\
        );

    \I__11719\ : CascadeMux
    port map (
            O => \N__51496\,
            I => \N__51380\
        );

    \I__11718\ : CascadeMux
    port map (
            O => \N__51495\,
            I => \N__51377\
        );

    \I__11717\ : InMux
    port map (
            O => \N__51494\,
            I => \N__51366\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__51489\,
            I => \N__51361\
        );

    \I__11715\ : LocalMux
    port map (
            O => \N__51486\,
            I => \N__51361\
        );

    \I__11714\ : Span4Mux_v
    port map (
            O => \N__51479\,
            I => \N__51352\
        );

    \I__11713\ : Span4Mux_h
    port map (
            O => \N__51476\,
            I => \N__51349\
        );

    \I__11712\ : InMux
    port map (
            O => \N__51475\,
            I => \N__51346\
        );

    \I__11711\ : CascadeMux
    port map (
            O => \N__51474\,
            I => \N__51335\
        );

    \I__11710\ : CascadeMux
    port map (
            O => \N__51473\,
            I => \N__51332\
        );

    \I__11709\ : CascadeMux
    port map (
            O => \N__51472\,
            I => \N__51329\
        );

    \I__11708\ : CascadeMux
    port map (
            O => \N__51471\,
            I => \N__51326\
        );

    \I__11707\ : CascadeMux
    port map (
            O => \N__51470\,
            I => \N__51323\
        );

    \I__11706\ : CascadeMux
    port map (
            O => \N__51469\,
            I => \N__51320\
        );

    \I__11705\ : CascadeMux
    port map (
            O => \N__51468\,
            I => \N__51317\
        );

    \I__11704\ : CascadeMux
    port map (
            O => \N__51467\,
            I => \N__51314\
        );

    \I__11703\ : CascadeMux
    port map (
            O => \N__51466\,
            I => \N__51311\
        );

    \I__11702\ : CascadeMux
    port map (
            O => \N__51465\,
            I => \N__51308\
        );

    \I__11701\ : CascadeMux
    port map (
            O => \N__51464\,
            I => \N__51305\
        );

    \I__11700\ : CascadeMux
    port map (
            O => \N__51463\,
            I => \N__51302\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__51454\,
            I => \N__51286\
        );

    \I__11698\ : Span4Mux_v
    port map (
            O => \N__51449\,
            I => \N__51277\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__51440\,
            I => \N__51277\
        );

    \I__11696\ : LocalMux
    port map (
            O => \N__51431\,
            I => \N__51277\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__51422\,
            I => \N__51277\
        );

    \I__11694\ : CascadeMux
    port map (
            O => \N__51421\,
            I => \N__51274\
        );

    \I__11693\ : CascadeMux
    port map (
            O => \N__51420\,
            I => \N__51271\
        );

    \I__11692\ : CascadeMux
    port map (
            O => \N__51419\,
            I => \N__51268\
        );

    \I__11691\ : CascadeMux
    port map (
            O => \N__51418\,
            I => \N__51265\
        );

    \I__11690\ : InMux
    port map (
            O => \N__51417\,
            I => \N__51250\
        );

    \I__11689\ : InMux
    port map (
            O => \N__51414\,
            I => \N__51250\
        );

    \I__11688\ : InMux
    port map (
            O => \N__51413\,
            I => \N__51250\
        );

    \I__11687\ : InMux
    port map (
            O => \N__51410\,
            I => \N__51250\
        );

    \I__11686\ : InMux
    port map (
            O => \N__51409\,
            I => \N__51250\
        );

    \I__11685\ : InMux
    port map (
            O => \N__51406\,
            I => \N__51250\
        );

    \I__11684\ : InMux
    port map (
            O => \N__51405\,
            I => \N__51250\
        );

    \I__11683\ : InMux
    port map (
            O => \N__51402\,
            I => \N__51233\
        );

    \I__11682\ : InMux
    port map (
            O => \N__51401\,
            I => \N__51233\
        );

    \I__11681\ : InMux
    port map (
            O => \N__51398\,
            I => \N__51233\
        );

    \I__11680\ : InMux
    port map (
            O => \N__51397\,
            I => \N__51233\
        );

    \I__11679\ : InMux
    port map (
            O => \N__51394\,
            I => \N__51233\
        );

    \I__11678\ : InMux
    port map (
            O => \N__51393\,
            I => \N__51233\
        );

    \I__11677\ : InMux
    port map (
            O => \N__51390\,
            I => \N__51233\
        );

    \I__11676\ : InMux
    port map (
            O => \N__51389\,
            I => \N__51233\
        );

    \I__11675\ : CascadeMux
    port map (
            O => \N__51388\,
            I => \N__51229\
        );

    \I__11674\ : CascadeMux
    port map (
            O => \N__51387\,
            I => \N__51225\
        );

    \I__11673\ : CascadeMux
    port map (
            O => \N__51386\,
            I => \N__51221\
        );

    \I__11672\ : InMux
    port map (
            O => \N__51383\,
            I => \N__51213\
        );

    \I__11671\ : InMux
    port map (
            O => \N__51380\,
            I => \N__51213\
        );

    \I__11670\ : InMux
    port map (
            O => \N__51377\,
            I => \N__51213\
        );

    \I__11669\ : CascadeMux
    port map (
            O => \N__51376\,
            I => \N__51210\
        );

    \I__11668\ : CascadeMux
    port map (
            O => \N__51375\,
            I => \N__51207\
        );

    \I__11667\ : CascadeMux
    port map (
            O => \N__51374\,
            I => \N__51204\
        );

    \I__11666\ : CascadeMux
    port map (
            O => \N__51373\,
            I => \N__51201\
        );

    \I__11665\ : InMux
    port map (
            O => \N__51372\,
            I => \N__51192\
        );

    \I__11664\ : InMux
    port map (
            O => \N__51371\,
            I => \N__51192\
        );

    \I__11663\ : InMux
    port map (
            O => \N__51370\,
            I => \N__51192\
        );

    \I__11662\ : InMux
    port map (
            O => \N__51369\,
            I => \N__51192\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__51366\,
            I => \N__51189\
        );

    \I__11660\ : Span4Mux_s1_h
    port map (
            O => \N__51361\,
            I => \N__51186\
        );

    \I__11659\ : InMux
    port map (
            O => \N__51360\,
            I => \N__51183\
        );

    \I__11658\ : InMux
    port map (
            O => \N__51359\,
            I => \N__51172\
        );

    \I__11657\ : InMux
    port map (
            O => \N__51358\,
            I => \N__51172\
        );

    \I__11656\ : InMux
    port map (
            O => \N__51357\,
            I => \N__51172\
        );

    \I__11655\ : InMux
    port map (
            O => \N__51356\,
            I => \N__51172\
        );

    \I__11654\ : InMux
    port map (
            O => \N__51355\,
            I => \N__51172\
        );

    \I__11653\ : Span4Mux_h
    port map (
            O => \N__51352\,
            I => \N__51161\
        );

    \I__11652\ : Span4Mux_v
    port map (
            O => \N__51349\,
            I => \N__51161\
        );

    \I__11651\ : LocalMux
    port map (
            O => \N__51346\,
            I => \N__51161\
        );

    \I__11650\ : InMux
    port map (
            O => \N__51345\,
            I => \N__51152\
        );

    \I__11649\ : InMux
    port map (
            O => \N__51344\,
            I => \N__51152\
        );

    \I__11648\ : InMux
    port map (
            O => \N__51343\,
            I => \N__51152\
        );

    \I__11647\ : InMux
    port map (
            O => \N__51342\,
            I => \N__51152\
        );

    \I__11646\ : InMux
    port map (
            O => \N__51341\,
            I => \N__51143\
        );

    \I__11645\ : InMux
    port map (
            O => \N__51340\,
            I => \N__51143\
        );

    \I__11644\ : InMux
    port map (
            O => \N__51339\,
            I => \N__51143\
        );

    \I__11643\ : InMux
    port map (
            O => \N__51338\,
            I => \N__51143\
        );

    \I__11642\ : InMux
    port map (
            O => \N__51335\,
            I => \N__51133\
        );

    \I__11641\ : InMux
    port map (
            O => \N__51332\,
            I => \N__51133\
        );

    \I__11640\ : InMux
    port map (
            O => \N__51329\,
            I => \N__51133\
        );

    \I__11639\ : InMux
    port map (
            O => \N__51326\,
            I => \N__51133\
        );

    \I__11638\ : InMux
    port map (
            O => \N__51323\,
            I => \N__51124\
        );

    \I__11637\ : InMux
    port map (
            O => \N__51320\,
            I => \N__51124\
        );

    \I__11636\ : InMux
    port map (
            O => \N__51317\,
            I => \N__51124\
        );

    \I__11635\ : InMux
    port map (
            O => \N__51314\,
            I => \N__51124\
        );

    \I__11634\ : InMux
    port map (
            O => \N__51311\,
            I => \N__51115\
        );

    \I__11633\ : InMux
    port map (
            O => \N__51308\,
            I => \N__51115\
        );

    \I__11632\ : InMux
    port map (
            O => \N__51305\,
            I => \N__51115\
        );

    \I__11631\ : InMux
    port map (
            O => \N__51302\,
            I => \N__51115\
        );

    \I__11630\ : CascadeMux
    port map (
            O => \N__51301\,
            I => \N__51112\
        );

    \I__11629\ : CascadeMux
    port map (
            O => \N__51300\,
            I => \N__51109\
        );

    \I__11628\ : CascadeMux
    port map (
            O => \N__51299\,
            I => \N__51106\
        );

    \I__11627\ : CascadeMux
    port map (
            O => \N__51298\,
            I => \N__51103\
        );

    \I__11626\ : CascadeMux
    port map (
            O => \N__51297\,
            I => \N__51100\
        );

    \I__11625\ : CascadeMux
    port map (
            O => \N__51296\,
            I => \N__51097\
        );

    \I__11624\ : CascadeMux
    port map (
            O => \N__51295\,
            I => \N__51094\
        );

    \I__11623\ : CascadeMux
    port map (
            O => \N__51294\,
            I => \N__51091\
        );

    \I__11622\ : InMux
    port map (
            O => \N__51293\,
            I => \N__51087\
        );

    \I__11621\ : InMux
    port map (
            O => \N__51292\,
            I => \N__51081\
        );

    \I__11620\ : CascadeMux
    port map (
            O => \N__51291\,
            I => \N__51071\
        );

    \I__11619\ : CascadeMux
    port map (
            O => \N__51290\,
            I => \N__51067\
        );

    \I__11618\ : CascadeMux
    port map (
            O => \N__51289\,
            I => \N__51063\
        );

    \I__11617\ : Span4Mux_v
    port map (
            O => \N__51286\,
            I => \N__51055\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__51277\,
            I => \N__51055\
        );

    \I__11615\ : InMux
    port map (
            O => \N__51274\,
            I => \N__51050\
        );

    \I__11614\ : InMux
    port map (
            O => \N__51271\,
            I => \N__51050\
        );

    \I__11613\ : InMux
    port map (
            O => \N__51268\,
            I => \N__51045\
        );

    \I__11612\ : InMux
    port map (
            O => \N__51265\,
            I => \N__51045\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__51250\,
            I => \N__51040\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__51233\,
            I => \N__51040\
        );

    \I__11609\ : InMux
    port map (
            O => \N__51232\,
            I => \N__51025\
        );

    \I__11608\ : InMux
    port map (
            O => \N__51229\,
            I => \N__51025\
        );

    \I__11607\ : InMux
    port map (
            O => \N__51228\,
            I => \N__51025\
        );

    \I__11606\ : InMux
    port map (
            O => \N__51225\,
            I => \N__51025\
        );

    \I__11605\ : InMux
    port map (
            O => \N__51224\,
            I => \N__51025\
        );

    \I__11604\ : InMux
    port map (
            O => \N__51221\,
            I => \N__51025\
        );

    \I__11603\ : InMux
    port map (
            O => \N__51220\,
            I => \N__51025\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__51213\,
            I => \N__51022\
        );

    \I__11601\ : InMux
    port map (
            O => \N__51210\,
            I => \N__51013\
        );

    \I__11600\ : InMux
    port map (
            O => \N__51207\,
            I => \N__51013\
        );

    \I__11599\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51013\
        );

    \I__11598\ : InMux
    port map (
            O => \N__51201\,
            I => \N__51013\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__51192\,
            I => \N__51010\
        );

    \I__11596\ : Span4Mux_v
    port map (
            O => \N__51189\,
            I => \N__51001\
        );

    \I__11595\ : Span4Mux_v
    port map (
            O => \N__51186\,
            I => \N__51001\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__51183\,
            I => \N__51001\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__51172\,
            I => \N__51001\
        );

    \I__11592\ : InMux
    port map (
            O => \N__51171\,
            I => \N__50998\
        );

    \I__11591\ : InMux
    port map (
            O => \N__51170\,
            I => \N__50993\
        );

    \I__11590\ : InMux
    port map (
            O => \N__51169\,
            I => \N__50993\
        );

    \I__11589\ : InMux
    port map (
            O => \N__51168\,
            I => \N__50990\
        );

    \I__11588\ : Span4Mux_h
    port map (
            O => \N__51161\,
            I => \N__50982\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__51152\,
            I => \N__50982\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__51143\,
            I => \N__50982\
        );

    \I__11585\ : InMux
    port map (
            O => \N__51142\,
            I => \N__50979\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__51133\,
            I => \N__50976\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__51124\,
            I => \N__50971\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__51115\,
            I => \N__50971\
        );

    \I__11581\ : InMux
    port map (
            O => \N__51112\,
            I => \N__50962\
        );

    \I__11580\ : InMux
    port map (
            O => \N__51109\,
            I => \N__50962\
        );

    \I__11579\ : InMux
    port map (
            O => \N__51106\,
            I => \N__50962\
        );

    \I__11578\ : InMux
    port map (
            O => \N__51103\,
            I => \N__50962\
        );

    \I__11577\ : InMux
    port map (
            O => \N__51100\,
            I => \N__50957\
        );

    \I__11576\ : InMux
    port map (
            O => \N__51097\,
            I => \N__50957\
        );

    \I__11575\ : InMux
    port map (
            O => \N__51094\,
            I => \N__50952\
        );

    \I__11574\ : InMux
    port map (
            O => \N__51091\,
            I => \N__50952\
        );

    \I__11573\ : InMux
    port map (
            O => \N__51090\,
            I => \N__50949\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__51087\,
            I => \N__50946\
        );

    \I__11571\ : InMux
    port map (
            O => \N__51086\,
            I => \N__50939\
        );

    \I__11570\ : InMux
    port map (
            O => \N__51085\,
            I => \N__50939\
        );

    \I__11569\ : InMux
    port map (
            O => \N__51084\,
            I => \N__50939\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__51081\,
            I => \N__50936\
        );

    \I__11567\ : InMux
    port map (
            O => \N__51080\,
            I => \N__50927\
        );

    \I__11566\ : InMux
    port map (
            O => \N__51079\,
            I => \N__50927\
        );

    \I__11565\ : InMux
    port map (
            O => \N__51078\,
            I => \N__50927\
        );

    \I__11564\ : InMux
    port map (
            O => \N__51077\,
            I => \N__50927\
        );

    \I__11563\ : InMux
    port map (
            O => \N__51076\,
            I => \N__50922\
        );

    \I__11562\ : InMux
    port map (
            O => \N__51075\,
            I => \N__50922\
        );

    \I__11561\ : InMux
    port map (
            O => \N__51074\,
            I => \N__50907\
        );

    \I__11560\ : InMux
    port map (
            O => \N__51071\,
            I => \N__50907\
        );

    \I__11559\ : InMux
    port map (
            O => \N__51070\,
            I => \N__50907\
        );

    \I__11558\ : InMux
    port map (
            O => \N__51067\,
            I => \N__50907\
        );

    \I__11557\ : InMux
    port map (
            O => \N__51066\,
            I => \N__50907\
        );

    \I__11556\ : InMux
    port map (
            O => \N__51063\,
            I => \N__50907\
        );

    \I__11555\ : InMux
    port map (
            O => \N__51062\,
            I => \N__50907\
        );

    \I__11554\ : CascadeMux
    port map (
            O => \N__51061\,
            I => \N__50904\
        );

    \I__11553\ : CascadeMux
    port map (
            O => \N__51060\,
            I => \N__50901\
        );

    \I__11552\ : Sp12to4
    port map (
            O => \N__51055\,
            I => \N__50893\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__51050\,
            I => \N__50893\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__51045\,
            I => \N__50893\
        );

    \I__11549\ : Span4Mux_v
    port map (
            O => \N__51040\,
            I => \N__50888\
        );

    \I__11548\ : LocalMux
    port map (
            O => \N__51025\,
            I => \N__50888\
        );

    \I__11547\ : Span4Mux_h
    port map (
            O => \N__51022\,
            I => \N__50885\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__51013\,
            I => \N__50882\
        );

    \I__11545\ : Span4Mux_v
    port map (
            O => \N__51010\,
            I => \N__50871\
        );

    \I__11544\ : Span4Mux_v
    port map (
            O => \N__51001\,
            I => \N__50871\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__50998\,
            I => \N__50871\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__50993\,
            I => \N__50871\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__50990\,
            I => \N__50871\
        );

    \I__11540\ : InMux
    port map (
            O => \N__50989\,
            I => \N__50868\
        );

    \I__11539\ : Span4Mux_h
    port map (
            O => \N__50982\,
            I => \N__50863\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__50979\,
            I => \N__50863\
        );

    \I__11537\ : Span4Mux_v
    port map (
            O => \N__50976\,
            I => \N__50852\
        );

    \I__11536\ : Span4Mux_h
    port map (
            O => \N__50971\,
            I => \N__50852\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__50962\,
            I => \N__50852\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__50957\,
            I => \N__50852\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__50952\,
            I => \N__50852\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__50949\,
            I => \N__50849\
        );

    \I__11531\ : Span4Mux_v
    port map (
            O => \N__50946\,
            I => \N__50844\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__50939\,
            I => \N__50844\
        );

    \I__11529\ : Span4Mux_v
    port map (
            O => \N__50936\,
            I => \N__50837\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__50927\,
            I => \N__50837\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__50922\,
            I => \N__50837\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__50907\,
            I => \N__50834\
        );

    \I__11525\ : InMux
    port map (
            O => \N__50904\,
            I => \N__50827\
        );

    \I__11524\ : InMux
    port map (
            O => \N__50901\,
            I => \N__50827\
        );

    \I__11523\ : InMux
    port map (
            O => \N__50900\,
            I => \N__50827\
        );

    \I__11522\ : Span12Mux_h
    port map (
            O => \N__50893\,
            I => \N__50824\
        );

    \I__11521\ : Span4Mux_v
    port map (
            O => \N__50888\,
            I => \N__50821\
        );

    \I__11520\ : Span4Mux_v
    port map (
            O => \N__50885\,
            I => \N__50818\
        );

    \I__11519\ : Span4Mux_v
    port map (
            O => \N__50882\,
            I => \N__50815\
        );

    \I__11518\ : Span4Mux_v
    port map (
            O => \N__50871\,
            I => \N__50810\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__50868\,
            I => \N__50810\
        );

    \I__11516\ : Span4Mux_h
    port map (
            O => \N__50863\,
            I => \N__50805\
        );

    \I__11515\ : Span4Mux_v
    port map (
            O => \N__50852\,
            I => \N__50805\
        );

    \I__11514\ : Span4Mux_v
    port map (
            O => \N__50849\,
            I => \N__50800\
        );

    \I__11513\ : Span4Mux_v
    port map (
            O => \N__50844\,
            I => \N__50800\
        );

    \I__11512\ : Span4Mux_v
    port map (
            O => \N__50837\,
            I => \N__50797\
        );

    \I__11511\ : Span4Mux_v
    port map (
            O => \N__50834\,
            I => \N__50794\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__50827\,
            I => \N__50791\
        );

    \I__11509\ : Span12Mux_v
    port map (
            O => \N__50824\,
            I => \N__50786\
        );

    \I__11508\ : Sp12to4
    port map (
            O => \N__50821\,
            I => \N__50786\
        );

    \I__11507\ : Span4Mux_v
    port map (
            O => \N__50818\,
            I => \N__50783\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__50815\,
            I => \N__50778\
        );

    \I__11505\ : Span4Mux_h
    port map (
            O => \N__50810\,
            I => \N__50778\
        );

    \I__11504\ : Span4Mux_v
    port map (
            O => \N__50805\,
            I => \N__50771\
        );

    \I__11503\ : Span4Mux_h
    port map (
            O => \N__50800\,
            I => \N__50771\
        );

    \I__11502\ : Span4Mux_h
    port map (
            O => \N__50797\,
            I => \N__50771\
        );

    \I__11501\ : Span4Mux_v
    port map (
            O => \N__50794\,
            I => \N__50766\
        );

    \I__11500\ : Span4Mux_v
    port map (
            O => \N__50791\,
            I => \N__50766\
        );

    \I__11499\ : Odrv12
    port map (
            O => \N__50786\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11498\ : Odrv4
    port map (
            O => \N__50783\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11497\ : Odrv4
    port map (
            O => \N__50778\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11496\ : Odrv4
    port map (
            O => \N__50771\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11495\ : Odrv4
    port map (
            O => \N__50766\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11494\ : InMux
    port map (
            O => \N__50755\,
            I => \N__50751\
        );

    \I__11493\ : InMux
    port map (
            O => \N__50754\,
            I => \N__50745\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__50751\,
            I => \N__50741\
        );

    \I__11491\ : InMux
    port map (
            O => \N__50750\,
            I => \N__50736\
        );

    \I__11490\ : InMux
    port map (
            O => \N__50749\,
            I => \N__50736\
        );

    \I__11489\ : InMux
    port map (
            O => \N__50748\,
            I => \N__50733\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__50745\,
            I => \N__50730\
        );

    \I__11487\ : InMux
    port map (
            O => \N__50744\,
            I => \N__50727\
        );

    \I__11486\ : Span4Mux_v
    port map (
            O => \N__50741\,
            I => \N__50722\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__50736\,
            I => \N__50722\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__50733\,
            I => \N__50719\
        );

    \I__11483\ : Span4Mux_h
    port map (
            O => \N__50730\,
            I => \N__50716\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__50727\,
            I => \N__50713\
        );

    \I__11481\ : Sp12to4
    port map (
            O => \N__50722\,
            I => \N__50708\
        );

    \I__11480\ : Span12Mux_s5_h
    port map (
            O => \N__50719\,
            I => \N__50708\
        );

    \I__11479\ : Span4Mux_v
    port map (
            O => \N__50716\,
            I => \N__50703\
        );

    \I__11478\ : Span4Mux_h
    port map (
            O => \N__50713\,
            I => \N__50703\
        );

    \I__11477\ : Odrv12
    port map (
            O => \N__50708\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__11476\ : Odrv4
    port map (
            O => \N__50703\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__11475\ : InMux
    port map (
            O => \N__50698\,
            I => \N__50695\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__50695\,
            I => \N__50691\
        );

    \I__11473\ : InMux
    port map (
            O => \N__50694\,
            I => \N__50688\
        );

    \I__11472\ : Span4Mux_v
    port map (
            O => \N__50691\,
            I => \N__50685\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__50688\,
            I => \N__50682\
        );

    \I__11470\ : Odrv4
    port map (
            O => \N__50685\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__11469\ : Odrv4
    port map (
            O => \N__50682\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__11468\ : CascadeMux
    port map (
            O => \N__50677\,
            I => \N__50673\
        );

    \I__11467\ : CascadeMux
    port map (
            O => \N__50676\,
            I => \N__50670\
        );

    \I__11466\ : InMux
    port map (
            O => \N__50673\,
            I => \N__50667\
        );

    \I__11465\ : InMux
    port map (
            O => \N__50670\,
            I => \N__50664\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__50667\,
            I => \N__50661\
        );

    \I__11463\ : LocalMux
    port map (
            O => \N__50664\,
            I => \N__50656\
        );

    \I__11462\ : Span4Mux_v
    port map (
            O => \N__50661\,
            I => \N__50656\
        );

    \I__11461\ : Span4Mux_h
    port map (
            O => \N__50656\,
            I => \N__50653\
        );

    \I__11460\ : Odrv4
    port map (
            O => \N__50653\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__11459\ : CascadeMux
    port map (
            O => \N__50650\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__11458\ : InMux
    port map (
            O => \N__50647\,
            I => \N__50638\
        );

    \I__11457\ : InMux
    port map (
            O => \N__50646\,
            I => \N__50638\
        );

    \I__11456\ : InMux
    port map (
            O => \N__50645\,
            I => \N__50638\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__50638\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__11454\ : InMux
    port map (
            O => \N__50635\,
            I => \N__50632\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__50632\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\
        );

    \I__11452\ : InMux
    port map (
            O => \N__50629\,
            I => \N__50626\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__50626\,
            I => \N__50623\
        );

    \I__11450\ : Odrv12
    port map (
            O => \N__50623\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\
        );

    \I__11449\ : InMux
    port map (
            O => \N__50620\,
            I => \N__50616\
        );

    \I__11448\ : InMux
    port map (
            O => \N__50619\,
            I => \N__50613\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__50616\,
            I => \N__50610\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__50613\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11445\ : Odrv4
    port map (
            O => \N__50610\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__11444\ : InMux
    port map (
            O => \N__50605\,
            I => \N__50602\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__50602\,
            I => \N__50599\
        );

    \I__11442\ : Odrv12
    port map (
            O => \N__50599\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\
        );

    \I__11441\ : InMux
    port map (
            O => \N__50596\,
            I => \N__50593\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__50593\,
            I => \N__50589\
        );

    \I__11439\ : CascadeMux
    port map (
            O => \N__50592\,
            I => \N__50586\
        );

    \I__11438\ : Span4Mux_h
    port map (
            O => \N__50589\,
            I => \N__50583\
        );

    \I__11437\ : InMux
    port map (
            O => \N__50586\,
            I => \N__50580\
        );

    \I__11436\ : Odrv4
    port map (
            O => \N__50583\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__50580\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__11434\ : InMux
    port map (
            O => \N__50575\,
            I => \N__50571\
        );

    \I__11433\ : InMux
    port map (
            O => \N__50574\,
            I => \N__50568\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__50571\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__50568\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__11430\ : InMux
    port map (
            O => \N__50563\,
            I => \N__50560\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__50560\,
            I => \N__50556\
        );

    \I__11428\ : InMux
    port map (
            O => \N__50559\,
            I => \N__50553\
        );

    \I__11427\ : Odrv4
    port map (
            O => \N__50556\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__50553\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__11425\ : InMux
    port map (
            O => \N__50548\,
            I => \N__50541\
        );

    \I__11424\ : InMux
    port map (
            O => \N__50547\,
            I => \N__50541\
        );

    \I__11423\ : CascadeMux
    port map (
            O => \N__50546\,
            I => \N__50533\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__50541\,
            I => \N__50519\
        );

    \I__11421\ : InMux
    port map (
            O => \N__50540\,
            I => \N__50510\
        );

    \I__11420\ : InMux
    port map (
            O => \N__50539\,
            I => \N__50510\
        );

    \I__11419\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50505\
        );

    \I__11418\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50505\
        );

    \I__11417\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50502\
        );

    \I__11416\ : InMux
    port map (
            O => \N__50533\,
            I => \N__50493\
        );

    \I__11415\ : InMux
    port map (
            O => \N__50532\,
            I => \N__50493\
        );

    \I__11414\ : InMux
    port map (
            O => \N__50531\,
            I => \N__50493\
        );

    \I__11413\ : InMux
    port map (
            O => \N__50530\,
            I => \N__50493\
        );

    \I__11412\ : InMux
    port map (
            O => \N__50529\,
            I => \N__50490\
        );

    \I__11411\ : CascadeMux
    port map (
            O => \N__50528\,
            I => \N__50487\
        );

    \I__11410\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50481\
        );

    \I__11409\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50474\
        );

    \I__11408\ : InMux
    port map (
            O => \N__50525\,
            I => \N__50469\
        );

    \I__11407\ : InMux
    port map (
            O => \N__50524\,
            I => \N__50469\
        );

    \I__11406\ : InMux
    port map (
            O => \N__50523\,
            I => \N__50464\
        );

    \I__11405\ : InMux
    port map (
            O => \N__50522\,
            I => \N__50464\
        );

    \I__11404\ : Span4Mux_h
    port map (
            O => \N__50519\,
            I => \N__50461\
        );

    \I__11403\ : InMux
    port map (
            O => \N__50518\,
            I => \N__50452\
        );

    \I__11402\ : InMux
    port map (
            O => \N__50517\,
            I => \N__50452\
        );

    \I__11401\ : InMux
    port map (
            O => \N__50516\,
            I => \N__50452\
        );

    \I__11400\ : InMux
    port map (
            O => \N__50515\,
            I => \N__50452\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__50510\,
            I => \N__50447\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__50505\,
            I => \N__50447\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__50502\,
            I => \N__50444\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__50493\,
            I => \N__50439\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__50490\,
            I => \N__50439\
        );

    \I__11394\ : InMux
    port map (
            O => \N__50487\,
            I => \N__50430\
        );

    \I__11393\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50430\
        );

    \I__11392\ : InMux
    port map (
            O => \N__50485\,
            I => \N__50430\
        );

    \I__11391\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50430\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__50481\,
            I => \N__50427\
        );

    \I__11389\ : InMux
    port map (
            O => \N__50480\,
            I => \N__50422\
        );

    \I__11388\ : InMux
    port map (
            O => \N__50479\,
            I => \N__50422\
        );

    \I__11387\ : InMux
    port map (
            O => \N__50478\,
            I => \N__50417\
        );

    \I__11386\ : InMux
    port map (
            O => \N__50477\,
            I => \N__50417\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__50474\,
            I => \N__50414\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__50469\,
            I => \N__50407\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__50464\,
            I => \N__50407\
        );

    \I__11382\ : Span4Mux_v
    port map (
            O => \N__50461\,
            I => \N__50407\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__50452\,
            I => \N__50398\
        );

    \I__11380\ : Span4Mux_v
    port map (
            O => \N__50447\,
            I => \N__50398\
        );

    \I__11379\ : Span4Mux_v
    port map (
            O => \N__50444\,
            I => \N__50398\
        );

    \I__11378\ : Span4Mux_h
    port map (
            O => \N__50439\,
            I => \N__50398\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__50430\,
            I => \N__50391\
        );

    \I__11376\ : Span12Mux_s10_v
    port map (
            O => \N__50427\,
            I => \N__50391\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__50422\,
            I => \N__50391\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__50417\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11373\ : Odrv4
    port map (
            O => \N__50414\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11372\ : Odrv4
    port map (
            O => \N__50407\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11371\ : Odrv4
    port map (
            O => \N__50398\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11370\ : Odrv12
    port map (
            O => \N__50391\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__11369\ : InMux
    port map (
            O => \N__50380\,
            I => \N__50376\
        );

    \I__11368\ : InMux
    port map (
            O => \N__50379\,
            I => \N__50373\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__50376\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__50373\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__11365\ : IoInMux
    port map (
            O => \N__50368\,
            I => \N__50365\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__50365\,
            I => \N__50362\
        );

    \I__11363\ : Span12Mux_s4_v
    port map (
            O => \N__50362\,
            I => \N__50359\
        );

    \I__11362\ : Span12Mux_v
    port map (
            O => \N__50359\,
            I => \N__50354\
        );

    \I__11361\ : InMux
    port map (
            O => \N__50358\,
            I => \N__50349\
        );

    \I__11360\ : InMux
    port map (
            O => \N__50357\,
            I => \N__50349\
        );

    \I__11359\ : Odrv12
    port map (
            O => \N__50354\,
            I => s1_phy_c
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__50349\,
            I => s1_phy_c
        );

    \I__11357\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50336\
        );

    \I__11356\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50336\
        );

    \I__11355\ : InMux
    port map (
            O => \N__50342\,
            I => \N__50333\
        );

    \I__11354\ : InMux
    port map (
            O => \N__50341\,
            I => \N__50329\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__50336\,
            I => \N__50323\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__50333\,
            I => \N__50323\
        );

    \I__11351\ : InMux
    port map (
            O => \N__50332\,
            I => \N__50320\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50317\
        );

    \I__11349\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50314\
        );

    \I__11348\ : Span12Mux_s6_h
    port map (
            O => \N__50323\,
            I => \N__50311\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__50320\,
            I => state_3
        );

    \I__11346\ : Odrv4
    port map (
            O => \N__50317\,
            I => state_3
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__50314\,
            I => state_3
        );

    \I__11344\ : Odrv12
    port map (
            O => \N__50311\,
            I => state_3
        );

    \I__11343\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50297\
        );

    \I__11342\ : CascadeMux
    port map (
            O => \N__50301\,
            I => \N__50293\
        );

    \I__11341\ : InMux
    port map (
            O => \N__50300\,
            I => \N__50290\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__50297\,
            I => \N__50287\
        );

    \I__11339\ : InMux
    port map (
            O => \N__50296\,
            I => \N__50282\
        );

    \I__11338\ : InMux
    port map (
            O => \N__50293\,
            I => \N__50282\
        );

    \I__11337\ : LocalMux
    port map (
            O => \N__50290\,
            I => \N__50279\
        );

    \I__11336\ : Span4Mux_h
    port map (
            O => \N__50287\,
            I => \N__50276\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__50282\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__11334\ : Odrv4
    port map (
            O => \N__50279\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__11333\ : Odrv4
    port map (
            O => \N__50276\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__11332\ : InMux
    port map (
            O => \N__50269\,
            I => \N__50263\
        );

    \I__11331\ : InMux
    port map (
            O => \N__50268\,
            I => \N__50256\
        );

    \I__11330\ : InMux
    port map (
            O => \N__50267\,
            I => \N__50256\
        );

    \I__11329\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50256\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__50263\,
            I => \N__50253\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__50256\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__11326\ : Odrv12
    port map (
            O => \N__50253\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__11325\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50245\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__50245\,
            I => \N__50240\
        );

    \I__11323\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50234\
        );

    \I__11322\ : InMux
    port map (
            O => \N__50243\,
            I => \N__50234\
        );

    \I__11321\ : Span4Mux_v
    port map (
            O => \N__50240\,
            I => \N__50231\
        );

    \I__11320\ : InMux
    port map (
            O => \N__50239\,
            I => \N__50228\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__50234\,
            I => \N__50223\
        );

    \I__11318\ : Span4Mux_v
    port map (
            O => \N__50231\,
            I => \N__50223\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__50228\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__11316\ : Odrv4
    port map (
            O => \N__50223\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__11315\ : InMux
    port map (
            O => \N__50218\,
            I => \N__50214\
        );

    \I__11314\ : InMux
    port map (
            O => \N__50217\,
            I => \N__50211\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__50214\,
            I => \N__50208\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__50211\,
            I => \N__50205\
        );

    \I__11311\ : Span12Mux_s10_h
    port map (
            O => \N__50208\,
            I => \N__50202\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__50205\,
            I => \N__50199\
        );

    \I__11309\ : Span12Mux_v
    port map (
            O => \N__50202\,
            I => \N__50196\
        );

    \I__11308\ : Odrv4
    port map (
            O => \N__50199\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__11307\ : Odrv12
    port map (
            O => \N__50196\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__11306\ : CascadeMux
    port map (
            O => \N__50191\,
            I => \N__50188\
        );

    \I__11305\ : InMux
    port map (
            O => \N__50188\,
            I => \N__50185\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__50185\,
            I => \N__50182\
        );

    \I__11303\ : Odrv4
    port map (
            O => \N__50182\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__11302\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50176\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__50176\,
            I => \N__50173\
        );

    \I__11300\ : Span4Mux_v
    port map (
            O => \N__50173\,
            I => \N__50170\
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__50170\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__11298\ : InMux
    port map (
            O => \N__50167\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__11297\ : InMux
    port map (
            O => \N__50164\,
            I => \N__50161\
        );

    \I__11296\ : LocalMux
    port map (
            O => \N__50161\,
            I => \N__50158\
        );

    \I__11295\ : Odrv4
    port map (
            O => \N__50158\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__11294\ : InMux
    port map (
            O => \N__50155\,
            I => \N__50152\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__50152\,
            I => \N__50149\
        );

    \I__11292\ : Span4Mux_v
    port map (
            O => \N__50149\,
            I => \N__50146\
        );

    \I__11291\ : Odrv4
    port map (
            O => \N__50146\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__11290\ : InMux
    port map (
            O => \N__50143\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__11289\ : CascadeMux
    port map (
            O => \N__50140\,
            I => \N__50137\
        );

    \I__11288\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50134\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__50134\,
            I => \N__50131\
        );

    \I__11286\ : Odrv4
    port map (
            O => \N__50131\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__11285\ : InMux
    port map (
            O => \N__50128\,
            I => \N__50125\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__50125\,
            I => \N__50122\
        );

    \I__11283\ : Span4Mux_h
    port map (
            O => \N__50122\,
            I => \N__50119\
        );

    \I__11282\ : Odrv4
    port map (
            O => \N__50119\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__11281\ : InMux
    port map (
            O => \N__50116\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__11280\ : CascadeMux
    port map (
            O => \N__50113\,
            I => \N__50109\
        );

    \I__11279\ : CascadeMux
    port map (
            O => \N__50112\,
            I => \N__50106\
        );

    \I__11278\ : InMux
    port map (
            O => \N__50109\,
            I => \N__50101\
        );

    \I__11277\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50097\
        );

    \I__11276\ : CascadeMux
    port map (
            O => \N__50105\,
            I => \N__50093\
        );

    \I__11275\ : CascadeMux
    port map (
            O => \N__50104\,
            I => \N__50070\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__50101\,
            I => \N__50063\
        );

    \I__11273\ : CascadeMux
    port map (
            O => \N__50100\,
            I => \N__50058\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__50097\,
            I => \N__50043\
        );

    \I__11271\ : InMux
    port map (
            O => \N__50096\,
            I => \N__50038\
        );

    \I__11270\ : InMux
    port map (
            O => \N__50093\,
            I => \N__50038\
        );

    \I__11269\ : CascadeMux
    port map (
            O => \N__50092\,
            I => \N__50034\
        );

    \I__11268\ : CascadeMux
    port map (
            O => \N__50091\,
            I => \N__50029\
        );

    \I__11267\ : CascadeMux
    port map (
            O => \N__50090\,
            I => \N__50026\
        );

    \I__11266\ : CascadeMux
    port map (
            O => \N__50089\,
            I => \N__50023\
        );

    \I__11265\ : CascadeMux
    port map (
            O => \N__50088\,
            I => \N__50020\
        );

    \I__11264\ : CascadeMux
    port map (
            O => \N__50087\,
            I => \N__50015\
        );

    \I__11263\ : CascadeMux
    port map (
            O => \N__50086\,
            I => \N__50008\
        );

    \I__11262\ : CascadeMux
    port map (
            O => \N__50085\,
            I => \N__49994\
        );

    \I__11261\ : InMux
    port map (
            O => \N__50084\,
            I => \N__49979\
        );

    \I__11260\ : InMux
    port map (
            O => \N__50083\,
            I => \N__49979\
        );

    \I__11259\ : InMux
    port map (
            O => \N__50082\,
            I => \N__49979\
        );

    \I__11258\ : InMux
    port map (
            O => \N__50081\,
            I => \N__49979\
        );

    \I__11257\ : InMux
    port map (
            O => \N__50080\,
            I => \N__49979\
        );

    \I__11256\ : InMux
    port map (
            O => \N__50079\,
            I => \N__49979\
        );

    \I__11255\ : InMux
    port map (
            O => \N__50078\,
            I => \N__49979\
        );

    \I__11254\ : InMux
    port map (
            O => \N__50077\,
            I => \N__49974\
        );

    \I__11253\ : InMux
    port map (
            O => \N__50076\,
            I => \N__49974\
        );

    \I__11252\ : InMux
    port map (
            O => \N__50075\,
            I => \N__49965\
        );

    \I__11251\ : InMux
    port map (
            O => \N__50074\,
            I => \N__49965\
        );

    \I__11250\ : InMux
    port map (
            O => \N__50073\,
            I => \N__49965\
        );

    \I__11249\ : InMux
    port map (
            O => \N__50070\,
            I => \N__49965\
        );

    \I__11248\ : CascadeMux
    port map (
            O => \N__50069\,
            I => \N__49960\
        );

    \I__11247\ : CascadeMux
    port map (
            O => \N__50068\,
            I => \N__49956\
        );

    \I__11246\ : CascadeMux
    port map (
            O => \N__50067\,
            I => \N__49952\
        );

    \I__11245\ : InMux
    port map (
            O => \N__50066\,
            I => \N__49944\
        );

    \I__11244\ : Span4Mux_v
    port map (
            O => \N__50063\,
            I => \N__49941\
        );

    \I__11243\ : InMux
    port map (
            O => \N__50062\,
            I => \N__49930\
        );

    \I__11242\ : InMux
    port map (
            O => \N__50061\,
            I => \N__49930\
        );

    \I__11241\ : InMux
    port map (
            O => \N__50058\,
            I => \N__49930\
        );

    \I__11240\ : InMux
    port map (
            O => \N__50057\,
            I => \N__49930\
        );

    \I__11239\ : InMux
    port map (
            O => \N__50056\,
            I => \N__49930\
        );

    \I__11238\ : InMux
    port map (
            O => \N__50055\,
            I => \N__49923\
        );

    \I__11237\ : InMux
    port map (
            O => \N__50054\,
            I => \N__49923\
        );

    \I__11236\ : InMux
    port map (
            O => \N__50053\,
            I => \N__49923\
        );

    \I__11235\ : CascadeMux
    port map (
            O => \N__50052\,
            I => \N__49919\
        );

    \I__11234\ : CascadeMux
    port map (
            O => \N__50051\,
            I => \N__49915\
        );

    \I__11233\ : CascadeMux
    port map (
            O => \N__50050\,
            I => \N__49911\
        );

    \I__11232\ : CascadeMux
    port map (
            O => \N__50049\,
            I => \N__49907\
        );

    \I__11231\ : CascadeMux
    port map (
            O => \N__50048\,
            I => \N__49903\
        );

    \I__11230\ : CascadeMux
    port map (
            O => \N__50047\,
            I => \N__49899\
        );

    \I__11229\ : CascadeMux
    port map (
            O => \N__50046\,
            I => \N__49895\
        );

    \I__11228\ : Span4Mux_v
    port map (
            O => \N__50043\,
            I => \N__49878\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__50038\,
            I => \N__49874\
        );

    \I__11226\ : InMux
    port map (
            O => \N__50037\,
            I => \N__49861\
        );

    \I__11225\ : InMux
    port map (
            O => \N__50034\,
            I => \N__49861\
        );

    \I__11224\ : InMux
    port map (
            O => \N__50033\,
            I => \N__49861\
        );

    \I__11223\ : InMux
    port map (
            O => \N__50032\,
            I => \N__49861\
        );

    \I__11222\ : InMux
    port map (
            O => \N__50029\,
            I => \N__49861\
        );

    \I__11221\ : InMux
    port map (
            O => \N__50026\,
            I => \N__49861\
        );

    \I__11220\ : InMux
    port map (
            O => \N__50023\,
            I => \N__49850\
        );

    \I__11219\ : InMux
    port map (
            O => \N__50020\,
            I => \N__49850\
        );

    \I__11218\ : InMux
    port map (
            O => \N__50019\,
            I => \N__49850\
        );

    \I__11217\ : InMux
    port map (
            O => \N__50018\,
            I => \N__49850\
        );

    \I__11216\ : InMux
    port map (
            O => \N__50015\,
            I => \N__49850\
        );

    \I__11215\ : InMux
    port map (
            O => \N__50014\,
            I => \N__49833\
        );

    \I__11214\ : InMux
    port map (
            O => \N__50013\,
            I => \N__49833\
        );

    \I__11213\ : InMux
    port map (
            O => \N__50012\,
            I => \N__49833\
        );

    \I__11212\ : InMux
    port map (
            O => \N__50011\,
            I => \N__49833\
        );

    \I__11211\ : InMux
    port map (
            O => \N__50008\,
            I => \N__49833\
        );

    \I__11210\ : InMux
    port map (
            O => \N__50007\,
            I => \N__49833\
        );

    \I__11209\ : InMux
    port map (
            O => \N__50006\,
            I => \N__49833\
        );

    \I__11208\ : InMux
    port map (
            O => \N__50005\,
            I => \N__49833\
        );

    \I__11207\ : CascadeMux
    port map (
            O => \N__50004\,
            I => \N__49830\
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__50003\,
            I => \N__49826\
        );

    \I__11205\ : CascadeMux
    port map (
            O => \N__50002\,
            I => \N__49821\
        );

    \I__11204\ : CascadeMux
    port map (
            O => \N__50001\,
            I => \N__49818\
        );

    \I__11203\ : CascadeMux
    port map (
            O => \N__50000\,
            I => \N__49814\
        );

    \I__11202\ : InMux
    port map (
            O => \N__49999\,
            I => \N__49805\
        );

    \I__11201\ : InMux
    port map (
            O => \N__49998\,
            I => \N__49805\
        );

    \I__11200\ : InMux
    port map (
            O => \N__49997\,
            I => \N__49805\
        );

    \I__11199\ : InMux
    port map (
            O => \N__49994\,
            I => \N__49805\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__49979\,
            I => \N__49800\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__49974\,
            I => \N__49800\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__49965\,
            I => \N__49797\
        );

    \I__11195\ : InMux
    port map (
            O => \N__49964\,
            I => \N__49780\
        );

    \I__11194\ : InMux
    port map (
            O => \N__49963\,
            I => \N__49780\
        );

    \I__11193\ : InMux
    port map (
            O => \N__49960\,
            I => \N__49780\
        );

    \I__11192\ : InMux
    port map (
            O => \N__49959\,
            I => \N__49780\
        );

    \I__11191\ : InMux
    port map (
            O => \N__49956\,
            I => \N__49780\
        );

    \I__11190\ : InMux
    port map (
            O => \N__49955\,
            I => \N__49780\
        );

    \I__11189\ : InMux
    port map (
            O => \N__49952\,
            I => \N__49780\
        );

    \I__11188\ : InMux
    port map (
            O => \N__49951\,
            I => \N__49780\
        );

    \I__11187\ : CascadeMux
    port map (
            O => \N__49950\,
            I => \N__49776\
        );

    \I__11186\ : CascadeMux
    port map (
            O => \N__49949\,
            I => \N__49772\
        );

    \I__11185\ : CascadeMux
    port map (
            O => \N__49948\,
            I => \N__49768\
        );

    \I__11184\ : CascadeMux
    port map (
            O => \N__49947\,
            I => \N__49764\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__49944\,
            I => \N__49761\
        );

    \I__11182\ : Span4Mux_h
    port map (
            O => \N__49941\,
            I => \N__49754\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__49930\,
            I => \N__49754\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__49923\,
            I => \N__49754\
        );

    \I__11179\ : InMux
    port map (
            O => \N__49922\,
            I => \N__49739\
        );

    \I__11178\ : InMux
    port map (
            O => \N__49919\,
            I => \N__49739\
        );

    \I__11177\ : InMux
    port map (
            O => \N__49918\,
            I => \N__49739\
        );

    \I__11176\ : InMux
    port map (
            O => \N__49915\,
            I => \N__49739\
        );

    \I__11175\ : InMux
    port map (
            O => \N__49914\,
            I => \N__49739\
        );

    \I__11174\ : InMux
    port map (
            O => \N__49911\,
            I => \N__49739\
        );

    \I__11173\ : InMux
    port map (
            O => \N__49910\,
            I => \N__49739\
        );

    \I__11172\ : InMux
    port map (
            O => \N__49907\,
            I => \N__49722\
        );

    \I__11171\ : InMux
    port map (
            O => \N__49906\,
            I => \N__49722\
        );

    \I__11170\ : InMux
    port map (
            O => \N__49903\,
            I => \N__49722\
        );

    \I__11169\ : InMux
    port map (
            O => \N__49902\,
            I => \N__49722\
        );

    \I__11168\ : InMux
    port map (
            O => \N__49899\,
            I => \N__49722\
        );

    \I__11167\ : InMux
    port map (
            O => \N__49898\,
            I => \N__49722\
        );

    \I__11166\ : InMux
    port map (
            O => \N__49895\,
            I => \N__49722\
        );

    \I__11165\ : InMux
    port map (
            O => \N__49894\,
            I => \N__49722\
        );

    \I__11164\ : CascadeMux
    port map (
            O => \N__49893\,
            I => \N__49719\
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__49892\,
            I => \N__49715\
        );

    \I__11162\ : CascadeMux
    port map (
            O => \N__49891\,
            I => \N__49711\
        );

    \I__11161\ : CascadeMux
    port map (
            O => \N__49890\,
            I => \N__49707\
        );

    \I__11160\ : CascadeMux
    port map (
            O => \N__49889\,
            I => \N__49703\
        );

    \I__11159\ : CascadeMux
    port map (
            O => \N__49888\,
            I => \N__49699\
        );

    \I__11158\ : CascadeMux
    port map (
            O => \N__49887\,
            I => \N__49695\
        );

    \I__11157\ : CascadeMux
    port map (
            O => \N__49886\,
            I => \N__49691\
        );

    \I__11156\ : CascadeMux
    port map (
            O => \N__49885\,
            I => \N__49685\
        );

    \I__11155\ : CascadeMux
    port map (
            O => \N__49884\,
            I => \N__49681\
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__49883\,
            I => \N__49676\
        );

    \I__11153\ : CascadeMux
    port map (
            O => \N__49882\,
            I => \N__49672\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__49881\,
            I => \N__49668\
        );

    \I__11151\ : Span4Mux_v
    port map (
            O => \N__49878\,
            I => \N__49665\
        );

    \I__11150\ : InMux
    port map (
            O => \N__49877\,
            I => \N__49662\
        );

    \I__11149\ : Span4Mux_v
    port map (
            O => \N__49874\,
            I => \N__49653\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__49861\,
            I => \N__49653\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__49850\,
            I => \N__49653\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__49833\,
            I => \N__49653\
        );

    \I__11145\ : InMux
    port map (
            O => \N__49830\,
            I => \N__49650\
        );

    \I__11144\ : InMux
    port map (
            O => \N__49829\,
            I => \N__49633\
        );

    \I__11143\ : InMux
    port map (
            O => \N__49826\,
            I => \N__49633\
        );

    \I__11142\ : InMux
    port map (
            O => \N__49825\,
            I => \N__49633\
        );

    \I__11141\ : InMux
    port map (
            O => \N__49824\,
            I => \N__49633\
        );

    \I__11140\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49633\
        );

    \I__11139\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49633\
        );

    \I__11138\ : InMux
    port map (
            O => \N__49817\,
            I => \N__49633\
        );

    \I__11137\ : InMux
    port map (
            O => \N__49814\,
            I => \N__49633\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__49805\,
            I => \N__49628\
        );

    \I__11135\ : Span4Mux_v
    port map (
            O => \N__49800\,
            I => \N__49628\
        );

    \I__11134\ : Span4Mux_v
    port map (
            O => \N__49797\,
            I => \N__49623\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__49780\,
            I => \N__49623\
        );

    \I__11132\ : InMux
    port map (
            O => \N__49779\,
            I => \N__49606\
        );

    \I__11131\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49606\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49606\
        );

    \I__11129\ : InMux
    port map (
            O => \N__49772\,
            I => \N__49606\
        );

    \I__11128\ : InMux
    port map (
            O => \N__49771\,
            I => \N__49606\
        );

    \I__11127\ : InMux
    port map (
            O => \N__49768\,
            I => \N__49606\
        );

    \I__11126\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49606\
        );

    \I__11125\ : InMux
    port map (
            O => \N__49764\,
            I => \N__49606\
        );

    \I__11124\ : Sp12to4
    port map (
            O => \N__49761\,
            I => \N__49597\
        );

    \I__11123\ : Sp12to4
    port map (
            O => \N__49754\,
            I => \N__49597\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__49739\,
            I => \N__49597\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__49722\,
            I => \N__49597\
        );

    \I__11120\ : InMux
    port map (
            O => \N__49719\,
            I => \N__49580\
        );

    \I__11119\ : InMux
    port map (
            O => \N__49718\,
            I => \N__49580\
        );

    \I__11118\ : InMux
    port map (
            O => \N__49715\,
            I => \N__49580\
        );

    \I__11117\ : InMux
    port map (
            O => \N__49714\,
            I => \N__49580\
        );

    \I__11116\ : InMux
    port map (
            O => \N__49711\,
            I => \N__49580\
        );

    \I__11115\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49580\
        );

    \I__11114\ : InMux
    port map (
            O => \N__49707\,
            I => \N__49580\
        );

    \I__11113\ : InMux
    port map (
            O => \N__49706\,
            I => \N__49580\
        );

    \I__11112\ : InMux
    port map (
            O => \N__49703\,
            I => \N__49563\
        );

    \I__11111\ : InMux
    port map (
            O => \N__49702\,
            I => \N__49563\
        );

    \I__11110\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49563\
        );

    \I__11109\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49563\
        );

    \I__11108\ : InMux
    port map (
            O => \N__49695\,
            I => \N__49563\
        );

    \I__11107\ : InMux
    port map (
            O => \N__49694\,
            I => \N__49563\
        );

    \I__11106\ : InMux
    port map (
            O => \N__49691\,
            I => \N__49563\
        );

    \I__11105\ : InMux
    port map (
            O => \N__49690\,
            I => \N__49563\
        );

    \I__11104\ : InMux
    port map (
            O => \N__49689\,
            I => \N__49560\
        );

    \I__11103\ : InMux
    port map (
            O => \N__49688\,
            I => \N__49549\
        );

    \I__11102\ : InMux
    port map (
            O => \N__49685\,
            I => \N__49549\
        );

    \I__11101\ : InMux
    port map (
            O => \N__49684\,
            I => \N__49549\
        );

    \I__11100\ : InMux
    port map (
            O => \N__49681\,
            I => \N__49549\
        );

    \I__11099\ : InMux
    port map (
            O => \N__49680\,
            I => \N__49549\
        );

    \I__11098\ : InMux
    port map (
            O => \N__49679\,
            I => \N__49536\
        );

    \I__11097\ : InMux
    port map (
            O => \N__49676\,
            I => \N__49536\
        );

    \I__11096\ : InMux
    port map (
            O => \N__49675\,
            I => \N__49536\
        );

    \I__11095\ : InMux
    port map (
            O => \N__49672\,
            I => \N__49536\
        );

    \I__11094\ : InMux
    port map (
            O => \N__49671\,
            I => \N__49536\
        );

    \I__11093\ : InMux
    port map (
            O => \N__49668\,
            I => \N__49536\
        );

    \I__11092\ : Odrv4
    port map (
            O => \N__49665\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__49662\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11090\ : Odrv4
    port map (
            O => \N__49653\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__49650\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__49633\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11087\ : Odrv4
    port map (
            O => \N__49628\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__49623\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__49606\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11084\ : Odrv12
    port map (
            O => \N__49597\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__49580\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__49563\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__49560\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__49549\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__49536\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11078\ : InMux
    port map (
            O => \N__49507\,
            I => \N__49483\
        );

    \I__11077\ : InMux
    port map (
            O => \N__49506\,
            I => \N__49483\
        );

    \I__11076\ : InMux
    port map (
            O => \N__49505\,
            I => \N__49483\
        );

    \I__11075\ : InMux
    port map (
            O => \N__49504\,
            I => \N__49483\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49503\,
            I => \N__49483\
        );

    \I__11073\ : InMux
    port map (
            O => \N__49502\,
            I => \N__49480\
        );

    \I__11072\ : InMux
    port map (
            O => \N__49501\,
            I => \N__49473\
        );

    \I__11071\ : InMux
    port map (
            O => \N__49500\,
            I => \N__49473\
        );

    \I__11070\ : InMux
    port map (
            O => \N__49499\,
            I => \N__49473\
        );

    \I__11069\ : InMux
    port map (
            O => \N__49498\,
            I => \N__49460\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49497\,
            I => \N__49460\
        );

    \I__11067\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49457\
        );

    \I__11066\ : InMux
    port map (
            O => \N__49495\,
            I => \N__49454\
        );

    \I__11065\ : InMux
    port map (
            O => \N__49494\,
            I => \N__49449\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__49483\,
            I => \N__49439\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__49480\,
            I => \N__49439\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__49473\,
            I => \N__49439\
        );

    \I__11061\ : InMux
    port map (
            O => \N__49472\,
            I => \N__49422\
        );

    \I__11060\ : InMux
    port map (
            O => \N__49471\,
            I => \N__49422\
        );

    \I__11059\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49422\
        );

    \I__11058\ : InMux
    port map (
            O => \N__49469\,
            I => \N__49422\
        );

    \I__11057\ : InMux
    port map (
            O => \N__49468\,
            I => \N__49422\
        );

    \I__11056\ : InMux
    port map (
            O => \N__49467\,
            I => \N__49422\
        );

    \I__11055\ : InMux
    port map (
            O => \N__49466\,
            I => \N__49422\
        );

    \I__11054\ : InMux
    port map (
            O => \N__49465\,
            I => \N__49422\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__49460\,
            I => \N__49419\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__49457\,
            I => \N__49416\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__49454\,
            I => \N__49405\
        );

    \I__11050\ : InMux
    port map (
            O => \N__49453\,
            I => \N__49400\
        );

    \I__11049\ : InMux
    port map (
            O => \N__49452\,
            I => \N__49400\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__49449\,
            I => \N__49397\
        );

    \I__11047\ : InMux
    port map (
            O => \N__49448\,
            I => \N__49390\
        );

    \I__11046\ : InMux
    port map (
            O => \N__49447\,
            I => \N__49390\
        );

    \I__11045\ : InMux
    port map (
            O => \N__49446\,
            I => \N__49390\
        );

    \I__11044\ : Span4Mux_v
    port map (
            O => \N__49439\,
            I => \N__49381\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__49422\,
            I => \N__49381\
        );

    \I__11042\ : Span4Mux_v
    port map (
            O => \N__49419\,
            I => \N__49381\
        );

    \I__11041\ : Span4Mux_h
    port map (
            O => \N__49416\,
            I => \N__49381\
        );

    \I__11040\ : InMux
    port map (
            O => \N__49415\,
            I => \N__49355\
        );

    \I__11039\ : InMux
    port map (
            O => \N__49414\,
            I => \N__49355\
        );

    \I__11038\ : InMux
    port map (
            O => \N__49413\,
            I => \N__49334\
        );

    \I__11037\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49334\
        );

    \I__11036\ : InMux
    port map (
            O => \N__49411\,
            I => \N__49334\
        );

    \I__11035\ : InMux
    port map (
            O => \N__49410\,
            I => \N__49334\
        );

    \I__11034\ : InMux
    port map (
            O => \N__49409\,
            I => \N__49334\
        );

    \I__11033\ : CascadeMux
    port map (
            O => \N__49408\,
            I => \N__49328\
        );

    \I__11032\ : Span4Mux_h
    port map (
            O => \N__49405\,
            I => \N__49321\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__49400\,
            I => \N__49321\
        );

    \I__11030\ : Span4Mux_v
    port map (
            O => \N__49397\,
            I => \N__49316\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__49390\,
            I => \N__49316\
        );

    \I__11028\ : Span4Mux_v
    port map (
            O => \N__49381\,
            I => \N__49313\
        );

    \I__11027\ : InMux
    port map (
            O => \N__49380\,
            I => \N__49304\
        );

    \I__11026\ : InMux
    port map (
            O => \N__49379\,
            I => \N__49304\
        );

    \I__11025\ : InMux
    port map (
            O => \N__49378\,
            I => \N__49304\
        );

    \I__11024\ : InMux
    port map (
            O => \N__49377\,
            I => \N__49304\
        );

    \I__11023\ : InMux
    port map (
            O => \N__49376\,
            I => \N__49291\
        );

    \I__11022\ : InMux
    port map (
            O => \N__49375\,
            I => \N__49291\
        );

    \I__11021\ : InMux
    port map (
            O => \N__49374\,
            I => \N__49291\
        );

    \I__11020\ : InMux
    port map (
            O => \N__49373\,
            I => \N__49291\
        );

    \I__11019\ : InMux
    port map (
            O => \N__49372\,
            I => \N__49291\
        );

    \I__11018\ : InMux
    port map (
            O => \N__49371\,
            I => \N__49291\
        );

    \I__11017\ : InMux
    port map (
            O => \N__49370\,
            I => \N__49274\
        );

    \I__11016\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49274\
        );

    \I__11015\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49274\
        );

    \I__11014\ : InMux
    port map (
            O => \N__49367\,
            I => \N__49274\
        );

    \I__11013\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49274\
        );

    \I__11012\ : InMux
    port map (
            O => \N__49365\,
            I => \N__49274\
        );

    \I__11011\ : InMux
    port map (
            O => \N__49364\,
            I => \N__49274\
        );

    \I__11010\ : InMux
    port map (
            O => \N__49363\,
            I => \N__49274\
        );

    \I__11009\ : InMux
    port map (
            O => \N__49362\,
            I => \N__49267\
        );

    \I__11008\ : InMux
    port map (
            O => \N__49361\,
            I => \N__49267\
        );

    \I__11007\ : InMux
    port map (
            O => \N__49360\,
            I => \N__49267\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__49355\,
            I => \N__49264\
        );

    \I__11005\ : InMux
    port map (
            O => \N__49354\,
            I => \N__49249\
        );

    \I__11004\ : InMux
    port map (
            O => \N__49353\,
            I => \N__49249\
        );

    \I__11003\ : InMux
    port map (
            O => \N__49352\,
            I => \N__49249\
        );

    \I__11002\ : InMux
    port map (
            O => \N__49351\,
            I => \N__49249\
        );

    \I__11001\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49249\
        );

    \I__11000\ : InMux
    port map (
            O => \N__49349\,
            I => \N__49249\
        );

    \I__10999\ : InMux
    port map (
            O => \N__49348\,
            I => \N__49249\
        );

    \I__10998\ : InMux
    port map (
            O => \N__49347\,
            I => \N__49242\
        );

    \I__10997\ : InMux
    port map (
            O => \N__49346\,
            I => \N__49242\
        );

    \I__10996\ : InMux
    port map (
            O => \N__49345\,
            I => \N__49242\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__49334\,
            I => \N__49239\
        );

    \I__10994\ : InMux
    port map (
            O => \N__49333\,
            I => \N__49226\
        );

    \I__10993\ : InMux
    port map (
            O => \N__49332\,
            I => \N__49226\
        );

    \I__10992\ : InMux
    port map (
            O => \N__49331\,
            I => \N__49226\
        );

    \I__10991\ : InMux
    port map (
            O => \N__49328\,
            I => \N__49226\
        );

    \I__10990\ : InMux
    port map (
            O => \N__49327\,
            I => \N__49226\
        );

    \I__10989\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49226\
        );

    \I__10988\ : Span4Mux_v
    port map (
            O => \N__49321\,
            I => \N__49221\
        );

    \I__10987\ : Span4Mux_h
    port map (
            O => \N__49316\,
            I => \N__49221\
        );

    \I__10986\ : Odrv4
    port map (
            O => \N__49313\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__49304\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__49291\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__49274\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__49267\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10981\ : Odrv4
    port map (
            O => \N__49264\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__49249\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__49242\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10978\ : Odrv4
    port map (
            O => \N__49239\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__49226\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10976\ : Odrv4
    port map (
            O => \N__49221\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__10975\ : InMux
    port map (
            O => \N__49198\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__10974\ : InMux
    port map (
            O => \N__49195\,
            I => \N__49192\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__49192\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__10972\ : InMux
    port map (
            O => \N__49189\,
            I => \N__49186\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__49186\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__10970\ : InMux
    port map (
            O => \N__49183\,
            I => \N__49180\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__49180\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__10968\ : CascadeMux
    port map (
            O => \N__49177\,
            I => \N__49174\
        );

    \I__10967\ : InMux
    port map (
            O => \N__49174\,
            I => \N__49170\
        );

    \I__10966\ : InMux
    port map (
            O => \N__49173\,
            I => \N__49167\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__49170\,
            I => \N__49150\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__49167\,
            I => \N__49150\
        );

    \I__10963\ : InMux
    port map (
            O => \N__49166\,
            I => \N__49145\
        );

    \I__10962\ : InMux
    port map (
            O => \N__49165\,
            I => \N__49145\
        );

    \I__10961\ : InMux
    port map (
            O => \N__49164\,
            I => \N__49142\
        );

    \I__10960\ : InMux
    port map (
            O => \N__49163\,
            I => \N__49137\
        );

    \I__10959\ : InMux
    port map (
            O => \N__49162\,
            I => \N__49137\
        );

    \I__10958\ : InMux
    port map (
            O => \N__49161\,
            I => \N__49122\
        );

    \I__10957\ : InMux
    port map (
            O => \N__49160\,
            I => \N__49122\
        );

    \I__10956\ : InMux
    port map (
            O => \N__49159\,
            I => \N__49122\
        );

    \I__10955\ : InMux
    port map (
            O => \N__49158\,
            I => \N__49122\
        );

    \I__10954\ : InMux
    port map (
            O => \N__49157\,
            I => \N__49122\
        );

    \I__10953\ : InMux
    port map (
            O => \N__49156\,
            I => \N__49122\
        );

    \I__10952\ : InMux
    port map (
            O => \N__49155\,
            I => \N__49122\
        );

    \I__10951\ : Span4Mux_h
    port map (
            O => \N__49150\,
            I => \N__49101\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__49145\,
            I => \N__49098\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__49142\,
            I => \N__49091\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__49137\,
            I => \N__49091\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__49122\,
            I => \N__49091\
        );

    \I__10946\ : InMux
    port map (
            O => \N__49121\,
            I => \N__49080\
        );

    \I__10945\ : InMux
    port map (
            O => \N__49120\,
            I => \N__49080\
        );

    \I__10944\ : InMux
    port map (
            O => \N__49119\,
            I => \N__49080\
        );

    \I__10943\ : InMux
    port map (
            O => \N__49118\,
            I => \N__49080\
        );

    \I__10942\ : InMux
    port map (
            O => \N__49117\,
            I => \N__49080\
        );

    \I__10941\ : InMux
    port map (
            O => \N__49116\,
            I => \N__49063\
        );

    \I__10940\ : InMux
    port map (
            O => \N__49115\,
            I => \N__49063\
        );

    \I__10939\ : InMux
    port map (
            O => \N__49114\,
            I => \N__49063\
        );

    \I__10938\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49063\
        );

    \I__10937\ : InMux
    port map (
            O => \N__49112\,
            I => \N__49063\
        );

    \I__10936\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49063\
        );

    \I__10935\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49063\
        );

    \I__10934\ : InMux
    port map (
            O => \N__49109\,
            I => \N__49063\
        );

    \I__10933\ : InMux
    port map (
            O => \N__49108\,
            I => \N__49052\
        );

    \I__10932\ : InMux
    port map (
            O => \N__49107\,
            I => \N__49052\
        );

    \I__10931\ : InMux
    port map (
            O => \N__49106\,
            I => \N__49052\
        );

    \I__10930\ : InMux
    port map (
            O => \N__49105\,
            I => \N__49052\
        );

    \I__10929\ : InMux
    port map (
            O => \N__49104\,
            I => \N__49052\
        );

    \I__10928\ : Odrv4
    port map (
            O => \N__49101\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10927\ : Odrv4
    port map (
            O => \N__49098\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__49091\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10925\ : LocalMux
    port map (
            O => \N__49080\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__49063\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__49052\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__10922\ : InMux
    port map (
            O => \N__49039\,
            I => \N__49036\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__49036\,
            I => \N__49033\
        );

    \I__10920\ : Odrv12
    port map (
            O => \N__49033\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__10919\ : InMux
    port map (
            O => \N__49030\,
            I => \N__49027\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__49027\,
            I => \N__49024\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__49024\,
            I => \N__49020\
        );

    \I__10916\ : InMux
    port map (
            O => \N__49023\,
            I => \N__49017\
        );

    \I__10915\ : Odrv4
    port map (
            O => \N__49020\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__49017\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10913\ : InMux
    port map (
            O => \N__49012\,
            I => \N__49009\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__49009\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__10911\ : CascadeMux
    port map (
            O => \N__49006\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\
        );

    \I__10910\ : InMux
    port map (
            O => \N__49003\,
            I => \N__49000\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__49000\,
            I => \N__48997\
        );

    \I__10908\ : Odrv12
    port map (
            O => \N__48997\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\
        );

    \I__10907\ : InMux
    port map (
            O => \N__48994\,
            I => \N__48991\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__48991\,
            I => \N__48988\
        );

    \I__10905\ : Span12Mux_s9_v
    port map (
            O => \N__48988\,
            I => \N__48985\
        );

    \I__10904\ : Odrv12
    port map (
            O => \N__48985\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\
        );

    \I__10903\ : InMux
    port map (
            O => \N__48982\,
            I => \N__48979\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__48979\,
            I => \N__48976\
        );

    \I__10901\ : Span4Mux_h
    port map (
            O => \N__48976\,
            I => \N__48973\
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__48973\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__10899\ : InMux
    port map (
            O => \N__48970\,
            I => \N__48967\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__48967\,
            I => \N__48964\
        );

    \I__10897\ : Span4Mux_h
    port map (
            O => \N__48964\,
            I => \N__48961\
        );

    \I__10896\ : Odrv4
    port map (
            O => \N__48961\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__10895\ : InMux
    port map (
            O => \N__48958\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__10894\ : CascadeMux
    port map (
            O => \N__48955\,
            I => \N__48952\
        );

    \I__10893\ : InMux
    port map (
            O => \N__48952\,
            I => \N__48949\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__48949\,
            I => \N__48946\
        );

    \I__10891\ : Odrv4
    port map (
            O => \N__48946\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__10890\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48940\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__48940\,
            I => \N__48937\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__48937\,
            I => \N__48934\
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__48934\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__10886\ : InMux
    port map (
            O => \N__48931\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__10885\ : InMux
    port map (
            O => \N__48928\,
            I => \N__48925\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__48925\,
            I => \N__48922\
        );

    \I__10883\ : Odrv12
    port map (
            O => \N__48922\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__10882\ : InMux
    port map (
            O => \N__48919\,
            I => \N__48916\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__48916\,
            I => \N__48913\
        );

    \I__10880\ : Span4Mux_h
    port map (
            O => \N__48913\,
            I => \N__48910\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__48910\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__10878\ : InMux
    port map (
            O => \N__48907\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__10877\ : CascadeMux
    port map (
            O => \N__48904\,
            I => \N__48901\
        );

    \I__10876\ : InMux
    port map (
            O => \N__48901\,
            I => \N__48898\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__48898\,
            I => \N__48895\
        );

    \I__10874\ : Odrv12
    port map (
            O => \N__48895\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__10873\ : InMux
    port map (
            O => \N__48892\,
            I => \N__48889\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__48889\,
            I => \N__48886\
        );

    \I__10871\ : Span4Mux_h
    port map (
            O => \N__48886\,
            I => \N__48883\
        );

    \I__10870\ : Odrv4
    port map (
            O => \N__48883\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__10869\ : InMux
    port map (
            O => \N__48880\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__10868\ : CascadeMux
    port map (
            O => \N__48877\,
            I => \N__48874\
        );

    \I__10867\ : InMux
    port map (
            O => \N__48874\,
            I => \N__48871\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__48871\,
            I => \N__48868\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__48868\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__10864\ : InMux
    port map (
            O => \N__48865\,
            I => \N__48862\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__48862\,
            I => \N__48859\
        );

    \I__10862\ : Span4Mux_h
    port map (
            O => \N__48859\,
            I => \N__48856\
        );

    \I__10861\ : Odrv4
    port map (
            O => \N__48856\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__10860\ : InMux
    port map (
            O => \N__48853\,
            I => \bfn_18_20_0_\
        );

    \I__10859\ : InMux
    port map (
            O => \N__48850\,
            I => \N__48847\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__48847\,
            I => \N__48844\
        );

    \I__10857\ : Odrv4
    port map (
            O => \N__48844\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__10856\ : InMux
    port map (
            O => \N__48841\,
            I => \N__48838\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__48838\,
            I => \N__48835\
        );

    \I__10854\ : Span4Mux_h
    port map (
            O => \N__48835\,
            I => \N__48832\
        );

    \I__10853\ : Odrv4
    port map (
            O => \N__48832\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__10852\ : InMux
    port map (
            O => \N__48829\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__10851\ : CascadeMux
    port map (
            O => \N__48826\,
            I => \N__48823\
        );

    \I__10850\ : InMux
    port map (
            O => \N__48823\,
            I => \N__48820\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__48820\,
            I => \N__48817\
        );

    \I__10848\ : Odrv4
    port map (
            O => \N__48817\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__10847\ : InMux
    port map (
            O => \N__48814\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__10846\ : InMux
    port map (
            O => \N__48811\,
            I => \N__48808\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__48808\,
            I => \N__48805\
        );

    \I__10844\ : Span4Mux_v
    port map (
            O => \N__48805\,
            I => \N__48802\
        );

    \I__10843\ : Odrv4
    port map (
            O => \N__48802\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__10842\ : InMux
    port map (
            O => \N__48799\,
            I => \N__48796\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__48796\,
            I => \N__48793\
        );

    \I__10840\ : Odrv12
    port map (
            O => \N__48793\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__10839\ : InMux
    port map (
            O => \N__48790\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__10838\ : CascadeMux
    port map (
            O => \N__48787\,
            I => \N__48784\
        );

    \I__10837\ : InMux
    port map (
            O => \N__48784\,
            I => \N__48781\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48778\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__48778\,
            I => \N__48775\
        );

    \I__10834\ : Odrv4
    port map (
            O => \N__48775\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__10833\ : InMux
    port map (
            O => \N__48772\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__10832\ : InMux
    port map (
            O => \N__48769\,
            I => \N__48766\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__48766\,
            I => \N__48763\
        );

    \I__10830\ : Odrv4
    port map (
            O => \N__48763\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__10829\ : InMux
    port map (
            O => \N__48760\,
            I => \N__48757\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__48757\,
            I => \N__48754\
        );

    \I__10827\ : Span4Mux_v
    port map (
            O => \N__48754\,
            I => \N__48751\
        );

    \I__10826\ : Odrv4
    port map (
            O => \N__48751\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__10825\ : InMux
    port map (
            O => \N__48748\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__10824\ : CascadeMux
    port map (
            O => \N__48745\,
            I => \N__48742\
        );

    \I__10823\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48739\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48736\
        );

    \I__10821\ : Span4Mux_v
    port map (
            O => \N__48736\,
            I => \N__48733\
        );

    \I__10820\ : Odrv4
    port map (
            O => \N__48733\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__10819\ : InMux
    port map (
            O => \N__48730\,
            I => \N__48727\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__48727\,
            I => \N__48724\
        );

    \I__10817\ : Span4Mux_h
    port map (
            O => \N__48724\,
            I => \N__48721\
        );

    \I__10816\ : Odrv4
    port map (
            O => \N__48721\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__10815\ : InMux
    port map (
            O => \N__48718\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__10814\ : InMux
    port map (
            O => \N__48715\,
            I => \N__48712\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__48712\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__10812\ : InMux
    port map (
            O => \N__48709\,
            I => \N__48706\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__48706\,
            I => \N__48703\
        );

    \I__10810\ : Span4Mux_h
    port map (
            O => \N__48703\,
            I => \N__48700\
        );

    \I__10809\ : Odrv4
    port map (
            O => \N__48700\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__10808\ : InMux
    port map (
            O => \N__48697\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__10807\ : InMux
    port map (
            O => \N__48694\,
            I => \N__48691\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__48691\,
            I => \N__48688\
        );

    \I__10805\ : Odrv12
    port map (
            O => \N__48688\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__10804\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48682\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__48682\,
            I => \N__48679\
        );

    \I__10802\ : Span4Mux_h
    port map (
            O => \N__48679\,
            I => \N__48676\
        );

    \I__10801\ : Odrv4
    port map (
            O => \N__48676\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__10800\ : InMux
    port map (
            O => \N__48673\,
            I => \bfn_18_19_0_\
        );

    \I__10799\ : CascadeMux
    port map (
            O => \N__48670\,
            I => \N__48667\
        );

    \I__10798\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48664\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__48664\,
            I => \N__48661\
        );

    \I__10796\ : Odrv12
    port map (
            O => \N__48661\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__10795\ : InMux
    port map (
            O => \N__48658\,
            I => \N__48655\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__48655\,
            I => \N__48652\
        );

    \I__10793\ : Span4Mux_h
    port map (
            O => \N__48652\,
            I => \N__48649\
        );

    \I__10792\ : Odrv4
    port map (
            O => \N__48649\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__10791\ : InMux
    port map (
            O => \N__48646\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__10790\ : InMux
    port map (
            O => \N__48643\,
            I => \N__48640\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__48640\,
            I => \N__48637\
        );

    \I__10788\ : Odrv12
    port map (
            O => \N__48637\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__10787\ : InMux
    port map (
            O => \N__48634\,
            I => \N__48631\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__48631\,
            I => \N__48628\
        );

    \I__10785\ : Span4Mux_h
    port map (
            O => \N__48628\,
            I => \N__48625\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__48625\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__10783\ : InMux
    port map (
            O => \N__48622\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__10782\ : CascadeMux
    port map (
            O => \N__48619\,
            I => \N__48616\
        );

    \I__10781\ : InMux
    port map (
            O => \N__48616\,
            I => \N__48613\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__48613\,
            I => \N__48610\
        );

    \I__10779\ : Span4Mux_v
    port map (
            O => \N__48610\,
            I => \N__48607\
        );

    \I__10778\ : Odrv4
    port map (
            O => \N__48607\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__10777\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48601\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__48601\,
            I => \N__48598\
        );

    \I__10775\ : Span4Mux_v
    port map (
            O => \N__48598\,
            I => \N__48595\
        );

    \I__10774\ : Odrv4
    port map (
            O => \N__48595\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__10773\ : InMux
    port map (
            O => \N__48592\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__10772\ : CascadeMux
    port map (
            O => \N__48589\,
            I => \N__48586\
        );

    \I__10771\ : InMux
    port map (
            O => \N__48586\,
            I => \N__48583\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__48583\,
            I => \N__48580\
        );

    \I__10769\ : Odrv12
    port map (
            O => \N__48580\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__10768\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48574\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__48574\,
            I => \N__48571\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__48571\,
            I => \N__48568\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__48568\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__10764\ : InMux
    port map (
            O => \N__48565\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__10763\ : InMux
    port map (
            O => \N__48562\,
            I => \N__48559\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__48559\,
            I => \N__48556\
        );

    \I__10761\ : Odrv12
    port map (
            O => \N__48556\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__10760\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48550\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__48550\,
            I => \N__48547\
        );

    \I__10758\ : Span4Mux_v
    port map (
            O => \N__48547\,
            I => \N__48544\
        );

    \I__10757\ : Odrv4
    port map (
            O => \N__48544\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__10756\ : InMux
    port map (
            O => \N__48541\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__10755\ : CascadeMux
    port map (
            O => \N__48538\,
            I => \N__48535\
        );

    \I__10754\ : InMux
    port map (
            O => \N__48535\,
            I => \N__48532\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__48532\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__10752\ : InMux
    port map (
            O => \N__48529\,
            I => \N__48526\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__48526\,
            I => \N__48523\
        );

    \I__10750\ : Span4Mux_h
    port map (
            O => \N__48523\,
            I => \N__48520\
        );

    \I__10749\ : Odrv4
    port map (
            O => \N__48520\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__10748\ : InMux
    port map (
            O => \N__48517\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__10747\ : CascadeMux
    port map (
            O => \N__48514\,
            I => \N__48511\
        );

    \I__10746\ : InMux
    port map (
            O => \N__48511\,
            I => \N__48508\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__48508\,
            I => \N__48505\
        );

    \I__10744\ : Span4Mux_v
    port map (
            O => \N__48505\,
            I => \N__48502\
        );

    \I__10743\ : Odrv4
    port map (
            O => \N__48502\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__10742\ : InMux
    port map (
            O => \N__48499\,
            I => \N__48496\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__48496\,
            I => \N__48493\
        );

    \I__10740\ : Span4Mux_h
    port map (
            O => \N__48493\,
            I => \N__48490\
        );

    \I__10739\ : Odrv4
    port map (
            O => \N__48490\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__10738\ : InMux
    port map (
            O => \N__48487\,
            I => \bfn_18_18_0_\
        );

    \I__10737\ : InMux
    port map (
            O => \N__48484\,
            I => \N__48481\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__48481\,
            I => \N__48478\
        );

    \I__10735\ : Span4Mux_v
    port map (
            O => \N__48478\,
            I => \N__48475\
        );

    \I__10734\ : Odrv4
    port map (
            O => \N__48475\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48472\,
            I => \N__48469\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48466\
        );

    \I__10731\ : Span4Mux_h
    port map (
            O => \N__48466\,
            I => \N__48463\
        );

    \I__10730\ : Odrv4
    port map (
            O => \N__48463\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__10729\ : InMux
    port map (
            O => \N__48460\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__10728\ : CascadeMux
    port map (
            O => \N__48457\,
            I => \N__48454\
        );

    \I__10727\ : InMux
    port map (
            O => \N__48454\,
            I => \N__48451\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__48451\,
            I => \N__48448\
        );

    \I__10725\ : Odrv12
    port map (
            O => \N__48448\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__10724\ : InMux
    port map (
            O => \N__48445\,
            I => \N__48442\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__48442\,
            I => \N__48439\
        );

    \I__10722\ : Span4Mux_v
    port map (
            O => \N__48439\,
            I => \N__48436\
        );

    \I__10721\ : Odrv4
    port map (
            O => \N__48436\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__10720\ : InMux
    port map (
            O => \N__48433\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__10719\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48427\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__48427\,
            I => \N__48424\
        );

    \I__10717\ : Odrv12
    port map (
            O => \N__48424\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__10716\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48418\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__48418\,
            I => \N__48415\
        );

    \I__10714\ : Span4Mux_v
    port map (
            O => \N__48415\,
            I => \N__48412\
        );

    \I__10713\ : Odrv4
    port map (
            O => \N__48412\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__10712\ : InMux
    port map (
            O => \N__48409\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__10711\ : CascadeMux
    port map (
            O => \N__48406\,
            I => \N__48403\
        );

    \I__10710\ : InMux
    port map (
            O => \N__48403\,
            I => \N__48400\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__48400\,
            I => \N__48397\
        );

    \I__10708\ : Odrv4
    port map (
            O => \N__48397\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__10707\ : InMux
    port map (
            O => \N__48394\,
            I => \N__48390\
        );

    \I__10706\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48387\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__48390\,
            I => \N__48381\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__48387\,
            I => \N__48381\
        );

    \I__10703\ : InMux
    port map (
            O => \N__48386\,
            I => \N__48378\
        );

    \I__10702\ : Span4Mux_v
    port map (
            O => \N__48381\,
            I => \N__48373\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48373\
        );

    \I__10700\ : Span4Mux_h
    port map (
            O => \N__48373\,
            I => \N__48369\
        );

    \I__10699\ : InMux
    port map (
            O => \N__48372\,
            I => \N__48366\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__48369\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__48366\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__10696\ : InMux
    port map (
            O => \N__48361\,
            I => \N__48357\
        );

    \I__10695\ : CascadeMux
    port map (
            O => \N__48360\,
            I => \N__48354\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__48357\,
            I => \N__48351\
        );

    \I__10693\ : InMux
    port map (
            O => \N__48354\,
            I => \N__48347\
        );

    \I__10692\ : Span4Mux_h
    port map (
            O => \N__48351\,
            I => \N__48344\
        );

    \I__10691\ : InMux
    port map (
            O => \N__48350\,
            I => \N__48341\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__48347\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__10689\ : Odrv4
    port map (
            O => \N__48344\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__48341\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__10687\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48331\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__48331\,
            I => \N__48328\
        );

    \I__10685\ : Span4Mux_v
    port map (
            O => \N__48328\,
            I => \N__48323\
        );

    \I__10684\ : InMux
    port map (
            O => \N__48327\,
            I => \N__48318\
        );

    \I__10683\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48318\
        );

    \I__10682\ : Odrv4
    port map (
            O => \N__48323\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__48318\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__10680\ : CascadeMux
    port map (
            O => \N__48313\,
            I => \N__48310\
        );

    \I__10679\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48307\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__48307\,
            I => \N__48304\
        );

    \I__10677\ : Span4Mux_v
    port map (
            O => \N__48304\,
            I => \N__48298\
        );

    \I__10676\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48291\
        );

    \I__10675\ : InMux
    port map (
            O => \N__48302\,
            I => \N__48291\
        );

    \I__10674\ : InMux
    port map (
            O => \N__48301\,
            I => \N__48291\
        );

    \I__10673\ : Odrv4
    port map (
            O => \N__48298\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__48291\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__48286\,
            I => \N__48283\
        );

    \I__10670\ : InMux
    port map (
            O => \N__48283\,
            I => \N__48280\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__48280\,
            I => \N__48277\
        );

    \I__10668\ : Odrv4
    port map (
            O => \N__48277\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__10667\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48268\
        );

    \I__10666\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48268\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__48268\,
            I => \N__48265\
        );

    \I__10664\ : Span4Mux_h
    port map (
            O => \N__48265\,
            I => \N__48261\
        );

    \I__10663\ : InMux
    port map (
            O => \N__48264\,
            I => \N__48258\
        );

    \I__10662\ : Odrv4
    port map (
            O => \N__48261\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__48258\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__10660\ : CascadeMux
    port map (
            O => \N__48253\,
            I => \N__48250\
        );

    \I__10659\ : InMux
    port map (
            O => \N__48250\,
            I => \N__48244\
        );

    \I__10658\ : InMux
    port map (
            O => \N__48249\,
            I => \N__48244\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__48244\,
            I => \N__48239\
        );

    \I__10656\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48234\
        );

    \I__10655\ : InMux
    port map (
            O => \N__48242\,
            I => \N__48234\
        );

    \I__10654\ : Span4Mux_v
    port map (
            O => \N__48239\,
            I => \N__48231\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__48234\,
            I => \N__48228\
        );

    \I__10652\ : Odrv4
    port map (
            O => \N__48231\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__48228\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__10650\ : CascadeMux
    port map (
            O => \N__48223\,
            I => \N__48220\
        );

    \I__10649\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48217\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__48217\,
            I => \N__48214\
        );

    \I__10647\ : Span4Mux_v
    port map (
            O => \N__48214\,
            I => \N__48210\
        );

    \I__10646\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48207\
        );

    \I__10645\ : Span4Mux_v
    port map (
            O => \N__48210\,
            I => \N__48202\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__48207\,
            I => \N__48199\
        );

    \I__10643\ : InMux
    port map (
            O => \N__48206\,
            I => \N__48196\
        );

    \I__10642\ : InMux
    port map (
            O => \N__48205\,
            I => \N__48193\
        );

    \I__10641\ : Odrv4
    port map (
            O => \N__48202\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10640\ : Odrv4
    port map (
            O => \N__48199\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__48196\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__48193\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10637\ : CascadeMux
    port map (
            O => \N__48184\,
            I => \N__48181\
        );

    \I__10636\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48178\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__48178\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__10634\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48172\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__48172\,
            I => \N__48169\
        );

    \I__10632\ : Odrv4
    port map (
            O => \N__48169\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__48166\,
            I => \N__48163\
        );

    \I__10630\ : InMux
    port map (
            O => \N__48163\,
            I => \N__48160\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__48160\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__10628\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48154\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48151\
        );

    \I__10626\ : Span4Mux_v
    port map (
            O => \N__48151\,
            I => \N__48148\
        );

    \I__10625\ : Odrv4
    port map (
            O => \N__48148\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__10624\ : InMux
    port map (
            O => \N__48145\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__10623\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48139\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__48139\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__10621\ : InMux
    port map (
            O => \N__48136\,
            I => \N__48133\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__48133\,
            I => \N__48130\
        );

    \I__10619\ : Span4Mux_h
    port map (
            O => \N__48130\,
            I => \N__48127\
        );

    \I__10618\ : Odrv4
    port map (
            O => \N__48127\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__10617\ : InMux
    port map (
            O => \N__48124\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__10616\ : InMux
    port map (
            O => \N__48121\,
            I => \N__48118\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__48112\
        );

    \I__10614\ : InMux
    port map (
            O => \N__48117\,
            I => \N__48109\
        );

    \I__10613\ : InMux
    port map (
            O => \N__48116\,
            I => \N__48104\
        );

    \I__10612\ : InMux
    port map (
            O => \N__48115\,
            I => \N__48104\
        );

    \I__10611\ : Odrv12
    port map (
            O => \N__48112\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__48109\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__48104\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__10608\ : InMux
    port map (
            O => \N__48097\,
            I => \N__48093\
        );

    \I__10607\ : InMux
    port map (
            O => \N__48096\,
            I => \N__48090\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__48093\,
            I => \N__48087\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__48090\,
            I => \N__48084\
        );

    \I__10604\ : Span4Mux_h
    port map (
            O => \N__48087\,
            I => \N__48078\
        );

    \I__10603\ : Span4Mux_h
    port map (
            O => \N__48084\,
            I => \N__48078\
        );

    \I__10602\ : InMux
    port map (
            O => \N__48083\,
            I => \N__48075\
        );

    \I__10601\ : Odrv4
    port map (
            O => \N__48078\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__48075\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__10599\ : CascadeMux
    port map (
            O => \N__48070\,
            I => \N__48067\
        );

    \I__10598\ : InMux
    port map (
            O => \N__48067\,
            I => \N__48063\
        );

    \I__10597\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48060\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__48063\,
            I => \N__48054\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__48060\,
            I => \N__48054\
        );

    \I__10594\ : InMux
    port map (
            O => \N__48059\,
            I => \N__48051\
        );

    \I__10593\ : Span4Mux_v
    port map (
            O => \N__48054\,
            I => \N__48045\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__48051\,
            I => \N__48045\
        );

    \I__10591\ : InMux
    port map (
            O => \N__48050\,
            I => \N__48042\
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__48045\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__48042\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__48037\,
            I => \N__48034\
        );

    \I__10587\ : InMux
    port map (
            O => \N__48034\,
            I => \N__48029\
        );

    \I__10586\ : InMux
    port map (
            O => \N__48033\,
            I => \N__48026\
        );

    \I__10585\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48023\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__48029\,
            I => \N__48020\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__48026\,
            I => \N__48017\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__48023\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10581\ : Odrv12
    port map (
            O => \N__48020\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10580\ : Odrv4
    port map (
            O => \N__48017\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__10579\ : CascadeMux
    port map (
            O => \N__48010\,
            I => \N__48007\
        );

    \I__10578\ : InMux
    port map (
            O => \N__48007\,
            I => \N__48002\
        );

    \I__10577\ : InMux
    port map (
            O => \N__48006\,
            I => \N__47999\
        );

    \I__10576\ : InMux
    port map (
            O => \N__48005\,
            I => \N__47996\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__48002\,
            I => \N__47993\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__47999\,
            I => \N__47990\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__47996\,
            I => \N__47987\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__47993\,
            I => \N__47983\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__47990\,
            I => \N__47980\
        );

    \I__10570\ : Span4Mux_v
    port map (
            O => \N__47987\,
            I => \N__47977\
        );

    \I__10569\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47974\
        );

    \I__10568\ : Odrv4
    port map (
            O => \N__47983\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__47980\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10566\ : Odrv4
    port map (
            O => \N__47977\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__47974\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10564\ : InMux
    port map (
            O => \N__47965\,
            I => \N__47961\
        );

    \I__10563\ : InMux
    port map (
            O => \N__47964\,
            I => \N__47957\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__47961\,
            I => \N__47954\
        );

    \I__10561\ : InMux
    port map (
            O => \N__47960\,
            I => \N__47951\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__47957\,
            I => \N__47948\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__47954\,
            I => \N__47945\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__47951\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10557\ : Odrv4
    port map (
            O => \N__47948\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10556\ : Odrv4
    port map (
            O => \N__47945\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__10555\ : InMux
    port map (
            O => \N__47938\,
            I => \N__47935\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__47935\,
            I => \N__47931\
        );

    \I__10553\ : InMux
    port map (
            O => \N__47934\,
            I => \N__47927\
        );

    \I__10552\ : Span4Mux_v
    port map (
            O => \N__47931\,
            I => \N__47924\
        );

    \I__10551\ : InMux
    port map (
            O => \N__47930\,
            I => \N__47921\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__47927\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10549\ : Odrv4
    port map (
            O => \N__47924\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__47921\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__47914\,
            I => \N__47911\
        );

    \I__10546\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47907\
        );

    \I__10545\ : CascadeMux
    port map (
            O => \N__47910\,
            I => \N__47904\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__47907\,
            I => \N__47901\
        );

    \I__10543\ : InMux
    port map (
            O => \N__47904\,
            I => \N__47898\
        );

    \I__10542\ : Span4Mux_h
    port map (
            O => \N__47901\,
            I => \N__47894\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__47898\,
            I => \N__47891\
        );

    \I__10540\ : InMux
    port map (
            O => \N__47897\,
            I => \N__47888\
        );

    \I__10539\ : Span4Mux_h
    port map (
            O => \N__47894\,
            I => \N__47884\
        );

    \I__10538\ : Span4Mux_h
    port map (
            O => \N__47891\,
            I => \N__47879\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__47888\,
            I => \N__47879\
        );

    \I__10536\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47876\
        );

    \I__10535\ : Odrv4
    port map (
            O => \N__47884\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__47879\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__47876\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__10532\ : InMux
    port map (
            O => \N__47869\,
            I => \N__47862\
        );

    \I__10531\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47862\
        );

    \I__10530\ : InMux
    port map (
            O => \N__47867\,
            I => \N__47859\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__47862\,
            I => \N__47855\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__47859\,
            I => \N__47852\
        );

    \I__10527\ : InMux
    port map (
            O => \N__47858\,
            I => \N__47849\
        );

    \I__10526\ : Span4Mux_v
    port map (
            O => \N__47855\,
            I => \N__47846\
        );

    \I__10525\ : Span4Mux_v
    port map (
            O => \N__47852\,
            I => \N__47841\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__47849\,
            I => \N__47841\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__47846\,
            I => \N__47838\
        );

    \I__10522\ : Span4Mux_h
    port map (
            O => \N__47841\,
            I => \N__47835\
        );

    \I__10521\ : Odrv4
    port map (
            O => \N__47838\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__47835\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__10519\ : CascadeMux
    port map (
            O => \N__47830\,
            I => \N__47826\
        );

    \I__10518\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47822\
        );

    \I__10517\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47817\
        );

    \I__10516\ : InMux
    port map (
            O => \N__47825\,
            I => \N__47817\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__47822\,
            I => \N__47814\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__47817\,
            I => \N__47811\
        );

    \I__10513\ : Odrv4
    port map (
            O => \N__47814\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__47811\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__10511\ : InMux
    port map (
            O => \N__47806\,
            I => \N__47803\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__47803\,
            I => \N__47798\
        );

    \I__10509\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47795\
        );

    \I__10508\ : InMux
    port map (
            O => \N__47801\,
            I => \N__47792\
        );

    \I__10507\ : Span12Mux_s9_h
    port map (
            O => \N__47798\,
            I => \N__47789\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__47795\,
            I => \N__47786\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__47792\,
            I => \N__47783\
        );

    \I__10504\ : Odrv12
    port map (
            O => \N__47789\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10503\ : Odrv12
    port map (
            O => \N__47786\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10502\ : Odrv4
    port map (
            O => \N__47783\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__10501\ : CascadeMux
    port map (
            O => \N__47776\,
            I => \N__47772\
        );

    \I__10500\ : CascadeMux
    port map (
            O => \N__47775\,
            I => \N__47769\
        );

    \I__10499\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47765\
        );

    \I__10498\ : InMux
    port map (
            O => \N__47769\,
            I => \N__47762\
        );

    \I__10497\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47759\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__47765\,
            I => \N__47755\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__47762\,
            I => \N__47750\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47750\
        );

    \I__10493\ : InMux
    port map (
            O => \N__47758\,
            I => \N__47747\
        );

    \I__10492\ : Span4Mux_h
    port map (
            O => \N__47755\,
            I => \N__47744\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__47750\,
            I => \N__47741\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__47747\,
            I => \N__47738\
        );

    \I__10489\ : Odrv4
    port map (
            O => \N__47744\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10488\ : Odrv4
    port map (
            O => \N__47741\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__47738\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__10486\ : CascadeMux
    port map (
            O => \N__47731\,
            I => \N__47728\
        );

    \I__10485\ : InMux
    port map (
            O => \N__47728\,
            I => \N__47724\
        );

    \I__10484\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47721\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47716\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__47721\,
            I => \N__47713\
        );

    \I__10481\ : InMux
    port map (
            O => \N__47720\,
            I => \N__47710\
        );

    \I__10480\ : InMux
    port map (
            O => \N__47719\,
            I => \N__47707\
        );

    \I__10479\ : Odrv4
    port map (
            O => \N__47716\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10478\ : Odrv12
    port map (
            O => \N__47713\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__47710\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__47707\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__10475\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47695\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__47695\,
            I => \N__47691\
        );

    \I__10473\ : InMux
    port map (
            O => \N__47694\,
            I => \N__47688\
        );

    \I__10472\ : Span4Mux_h
    port map (
            O => \N__47691\,
            I => \N__47684\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__47688\,
            I => \N__47681\
        );

    \I__10470\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47678\
        );

    \I__10469\ : Odrv4
    port map (
            O => \N__47684\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10468\ : Odrv4
    port map (
            O => \N__47681\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__47678\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10466\ : CascadeMux
    port map (
            O => \N__47671\,
            I => \N__47668\
        );

    \I__10465\ : InMux
    port map (
            O => \N__47668\,
            I => \N__47665\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__47665\,
            I => \N__47661\
        );

    \I__10463\ : InMux
    port map (
            O => \N__47664\,
            I => \N__47657\
        );

    \I__10462\ : Span4Mux_h
    port map (
            O => \N__47661\,
            I => \N__47654\
        );

    \I__10461\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47651\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__47657\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10459\ : Odrv4
    port map (
            O => \N__47654\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__47651\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__10457\ : CascadeMux
    port map (
            O => \N__47644\,
            I => \N__47641\
        );

    \I__10456\ : InMux
    port map (
            O => \N__47641\,
            I => \N__47637\
        );

    \I__10455\ : InMux
    port map (
            O => \N__47640\,
            I => \N__47634\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47630\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__47634\,
            I => \N__47627\
        );

    \I__10452\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47624\
        );

    \I__10451\ : Span4Mux_h
    port map (
            O => \N__47630\,
            I => \N__47620\
        );

    \I__10450\ : Span4Mux_h
    port map (
            O => \N__47627\,
            I => \N__47615\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__47624\,
            I => \N__47615\
        );

    \I__10448\ : InMux
    port map (
            O => \N__47623\,
            I => \N__47612\
        );

    \I__10447\ : Odrv4
    port map (
            O => \N__47620\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10446\ : Odrv4
    port map (
            O => \N__47615\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__47612\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__10444\ : InMux
    port map (
            O => \N__47605\,
            I => \N__47601\
        );

    \I__10443\ : InMux
    port map (
            O => \N__47604\,
            I => \N__47598\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__47601\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__47598\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__10440\ : InMux
    port map (
            O => \N__47593\,
            I => \N__47590\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__47590\,
            I => \N__47587\
        );

    \I__10438\ : Span4Mux_h
    port map (
            O => \N__47587\,
            I => \N__47584\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__47584\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\
        );

    \I__10436\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47577\
        );

    \I__10435\ : InMux
    port map (
            O => \N__47580\,
            I => \N__47574\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__47577\,
            I => \N__47571\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__47574\,
            I => \N__47568\
        );

    \I__10432\ : Span4Mux_v
    port map (
            O => \N__47571\,
            I => \N__47565\
        );

    \I__10431\ : Span4Mux_v
    port map (
            O => \N__47568\,
            I => \N__47560\
        );

    \I__10430\ : Span4Mux_h
    port map (
            O => \N__47565\,
            I => \N__47557\
        );

    \I__10429\ : InMux
    port map (
            O => \N__47564\,
            I => \N__47552\
        );

    \I__10428\ : InMux
    port map (
            O => \N__47563\,
            I => \N__47552\
        );

    \I__10427\ : Span4Mux_v
    port map (
            O => \N__47560\,
            I => \N__47549\
        );

    \I__10426\ : Span4Mux_v
    port map (
            O => \N__47557\,
            I => \N__47546\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__47552\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__47549\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__47546\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__10422\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47536\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__47536\,
            I => \N__47531\
        );

    \I__10420\ : InMux
    port map (
            O => \N__47535\,
            I => \N__47528\
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__47534\,
            I => \N__47525\
        );

    \I__10418\ : Span4Mux_v
    port map (
            O => \N__47531\,
            I => \N__47519\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__47528\,
            I => \N__47519\
        );

    \I__10416\ : InMux
    port map (
            O => \N__47525\,
            I => \N__47514\
        );

    \I__10415\ : InMux
    port map (
            O => \N__47524\,
            I => \N__47514\
        );

    \I__10414\ : Span4Mux_h
    port map (
            O => \N__47519\,
            I => \N__47511\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__47514\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__47511\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__10411\ : InMux
    port map (
            O => \N__47506\,
            I => \N__47503\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__47503\,
            I => \N__47498\
        );

    \I__10409\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47493\
        );

    \I__10408\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47493\
        );

    \I__10407\ : Span4Mux_v
    port map (
            O => \N__47498\,
            I => \N__47490\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__47493\,
            I => \N__47487\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__47490\,
            I => \N__47484\
        );

    \I__10404\ : Span4Mux_v
    port map (
            O => \N__47487\,
            I => \N__47481\
        );

    \I__10403\ : Span4Mux_v
    port map (
            O => \N__47484\,
            I => \N__47478\
        );

    \I__10402\ : Span4Mux_v
    port map (
            O => \N__47481\,
            I => \N__47475\
        );

    \I__10401\ : Odrv4
    port map (
            O => \N__47478\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__47475\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__10399\ : CEMux
    port map (
            O => \N__47470\,
            I => \N__47464\
        );

    \I__10398\ : CEMux
    port map (
            O => \N__47469\,
            I => \N__47461\
        );

    \I__10397\ : CEMux
    port map (
            O => \N__47468\,
            I => \N__47458\
        );

    \I__10396\ : CEMux
    port map (
            O => \N__47467\,
            I => \N__47455\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__47464\,
            I => \N__47452\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__47461\,
            I => \N__47447\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__47458\,
            I => \N__47447\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__47455\,
            I => \N__47444\
        );

    \I__10391\ : Span4Mux_v
    port map (
            O => \N__47452\,
            I => \N__47437\
        );

    \I__10390\ : Span4Mux_v
    port map (
            O => \N__47447\,
            I => \N__47437\
        );

    \I__10389\ : Span4Mux_h
    port map (
            O => \N__47444\,
            I => \N__47437\
        );

    \I__10388\ : Odrv4
    port map (
            O => \N__47437\,
            I => \delay_measurement_inst.delay_hc_timer.N_166_i\
        );

    \I__10387\ : InMux
    port map (
            O => \N__47434\,
            I => \N__47430\
        );

    \I__10386\ : InMux
    port map (
            O => \N__47433\,
            I => \N__47427\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__47430\,
            I => \N__47421\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__47427\,
            I => \N__47421\
        );

    \I__10383\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47418\
        );

    \I__10382\ : Span4Mux_v
    port map (
            O => \N__47421\,
            I => \N__47413\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__47418\,
            I => \N__47413\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__47413\,
            I => \N__47409\
        );

    \I__10379\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47406\
        );

    \I__10378\ : Odrv4
    port map (
            O => \N__47409\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__47406\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__10376\ : CascadeMux
    port map (
            O => \N__47401\,
            I => \N__47397\
        );

    \I__10375\ : CascadeMux
    port map (
            O => \N__47400\,
            I => \N__47394\
        );

    \I__10374\ : InMux
    port map (
            O => \N__47397\,
            I => \N__47390\
        );

    \I__10373\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47387\
        );

    \I__10372\ : InMux
    port map (
            O => \N__47393\,
            I => \N__47384\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__47390\,
            I => \N__47379\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__47387\,
            I => \N__47379\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__47384\,
            I => \N__47376\
        );

    \I__10368\ : Odrv4
    port map (
            O => \N__47379\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10367\ : Odrv4
    port map (
            O => \N__47376\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__10366\ : CEMux
    port map (
            O => \N__47371\,
            I => \N__47368\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47364\
        );

    \I__10364\ : CEMux
    port map (
            O => \N__47367\,
            I => \N__47361\
        );

    \I__10363\ : Span4Mux_v
    port map (
            O => \N__47364\,
            I => \N__47357\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__47361\,
            I => \N__47354\
        );

    \I__10361\ : CEMux
    port map (
            O => \N__47360\,
            I => \N__47350\
        );

    \I__10360\ : Span4Mux_h
    port map (
            O => \N__47357\,
            I => \N__47345\
        );

    \I__10359\ : Span4Mux_h
    port map (
            O => \N__47354\,
            I => \N__47345\
        );

    \I__10358\ : CEMux
    port map (
            O => \N__47353\,
            I => \N__47342\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__47350\,
            I => \N__47339\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__47345\,
            I => \N__47336\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__47342\,
            I => \N__47333\
        );

    \I__10354\ : Span4Mux_h
    port map (
            O => \N__47339\,
            I => \N__47330\
        );

    \I__10353\ : Span4Mux_h
    port map (
            O => \N__47336\,
            I => \N__47327\
        );

    \I__10352\ : Odrv12
    port map (
            O => \N__47333\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10351\ : Odrv4
    port map (
            O => \N__47330\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10350\ : Odrv4
    port map (
            O => \N__47327\,
            I => \current_shift_inst.timer_s1.N_164_i\
        );

    \I__10349\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47316\
        );

    \I__10348\ : InMux
    port map (
            O => \N__47319\,
            I => \N__47312\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__47316\,
            I => \N__47309\
        );

    \I__10346\ : InMux
    port map (
            O => \N__47315\,
            I => \N__47306\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__47312\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10344\ : Odrv12
    port map (
            O => \N__47309\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__47306\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__10342\ : CascadeMux
    port map (
            O => \N__47299\,
            I => \N__47295\
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__47298\,
            I => \N__47292\
        );

    \I__10340\ : InMux
    port map (
            O => \N__47295\,
            I => \N__47289\
        );

    \I__10339\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47286\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__47289\,
            I => \N__47282\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__47286\,
            I => \N__47279\
        );

    \I__10336\ : InMux
    port map (
            O => \N__47285\,
            I => \N__47276\
        );

    \I__10335\ : Span4Mux_h
    port map (
            O => \N__47282\,
            I => \N__47270\
        );

    \I__10334\ : Span4Mux_h
    port map (
            O => \N__47279\,
            I => \N__47270\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__47276\,
            I => \N__47267\
        );

    \I__10332\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47264\
        );

    \I__10331\ : Odrv4
    port map (
            O => \N__47270\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10330\ : Odrv4
    port map (
            O => \N__47267\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__47264\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10328\ : InMux
    port map (
            O => \N__47257\,
            I => \N__47219\
        );

    \I__10327\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47219\
        );

    \I__10326\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47219\
        );

    \I__10325\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47219\
        );

    \I__10324\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47210\
        );

    \I__10323\ : InMux
    port map (
            O => \N__47252\,
            I => \N__47210\
        );

    \I__10322\ : InMux
    port map (
            O => \N__47251\,
            I => \N__47210\
        );

    \I__10321\ : InMux
    port map (
            O => \N__47250\,
            I => \N__47210\
        );

    \I__10320\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47201\
        );

    \I__10319\ : InMux
    port map (
            O => \N__47248\,
            I => \N__47201\
        );

    \I__10318\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47201\
        );

    \I__10317\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47201\
        );

    \I__10316\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47192\
        );

    \I__10315\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47192\
        );

    \I__10314\ : InMux
    port map (
            O => \N__47243\,
            I => \N__47192\
        );

    \I__10313\ : InMux
    port map (
            O => \N__47242\,
            I => \N__47192\
        );

    \I__10312\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47183\
        );

    \I__10311\ : InMux
    port map (
            O => \N__47240\,
            I => \N__47183\
        );

    \I__10310\ : InMux
    port map (
            O => \N__47239\,
            I => \N__47183\
        );

    \I__10309\ : InMux
    port map (
            O => \N__47238\,
            I => \N__47183\
        );

    \I__10308\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47174\
        );

    \I__10307\ : InMux
    port map (
            O => \N__47236\,
            I => \N__47174\
        );

    \I__10306\ : InMux
    port map (
            O => \N__47235\,
            I => \N__47174\
        );

    \I__10305\ : InMux
    port map (
            O => \N__47234\,
            I => \N__47174\
        );

    \I__10304\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47169\
        );

    \I__10303\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47169\
        );

    \I__10302\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47160\
        );

    \I__10301\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47160\
        );

    \I__10300\ : InMux
    port map (
            O => \N__47229\,
            I => \N__47160\
        );

    \I__10299\ : InMux
    port map (
            O => \N__47228\,
            I => \N__47160\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__47219\,
            I => \N__47157\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__47210\,
            I => \N__47146\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__47201\,
            I => \N__47146\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__47192\,
            I => \N__47146\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__47183\,
            I => \N__47146\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__47174\,
            I => \N__47146\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__47169\,
            I => \N__47137\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__47160\,
            I => \N__47137\
        );

    \I__10290\ : Span4Mux_v
    port map (
            O => \N__47157\,
            I => \N__47137\
        );

    \I__10289\ : Span4Mux_v
    port map (
            O => \N__47146\,
            I => \N__47137\
        );

    \I__10288\ : Span4Mux_h
    port map (
            O => \N__47137\,
            I => \N__47134\
        );

    \I__10287\ : Odrv4
    port map (
            O => \N__47134\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10286\ : InMux
    port map (
            O => \N__47131\,
            I => \N__47128\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__47128\,
            I => \N__47124\
        );

    \I__10284\ : InMux
    port map (
            O => \N__47127\,
            I => \N__47120\
        );

    \I__10283\ : Span4Mux_h
    port map (
            O => \N__47124\,
            I => \N__47117\
        );

    \I__10282\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47114\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__47120\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__47117\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__47114\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__10278\ : CascadeMux
    port map (
            O => \N__47107\,
            I => \N__47103\
        );

    \I__10277\ : CascadeMux
    port map (
            O => \N__47106\,
            I => \N__47100\
        );

    \I__10276\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47097\
        );

    \I__10275\ : InMux
    port map (
            O => \N__47100\,
            I => \N__47094\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__47097\,
            I => \N__47089\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__47094\,
            I => \N__47089\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__47089\,
            I => \N__47084\
        );

    \I__10271\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47079\
        );

    \I__10270\ : InMux
    port map (
            O => \N__47087\,
            I => \N__47079\
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__47084\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__47079\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__10267\ : CascadeMux
    port map (
            O => \N__47074\,
            I => \N__47071\
        );

    \I__10266\ : InMux
    port map (
            O => \N__47071\,
            I => \N__47067\
        );

    \I__10265\ : InMux
    port map (
            O => \N__47070\,
            I => \N__47064\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__47067\,
            I => \N__47058\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__47064\,
            I => \N__47058\
        );

    \I__10262\ : InMux
    port map (
            O => \N__47063\,
            I => \N__47055\
        );

    \I__10261\ : Span4Mux_h
    port map (
            O => \N__47058\,
            I => \N__47051\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__47048\
        );

    \I__10259\ : InMux
    port map (
            O => \N__47054\,
            I => \N__47045\
        );

    \I__10258\ : Odrv4
    port map (
            O => \N__47051\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10257\ : Odrv4
    port map (
            O => \N__47048\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__47045\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__10255\ : InMux
    port map (
            O => \N__47038\,
            I => \N__47033\
        );

    \I__10254\ : InMux
    port map (
            O => \N__47037\,
            I => \N__47030\
        );

    \I__10253\ : InMux
    port map (
            O => \N__47036\,
            I => \N__47027\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__47033\,
            I => \N__47022\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__47030\,
            I => \N__47022\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__47027\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__47022\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__10248\ : IoInMux
    port map (
            O => \N__47017\,
            I => \N__47014\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__47014\,
            I => \N__47011\
        );

    \I__10246\ : Span4Mux_s3_v
    port map (
            O => \N__47011\,
            I => \N__47008\
        );

    \I__10245\ : Sp12to4
    port map (
            O => \N__47008\,
            I => \N__47005\
        );

    \I__10244\ : Span12Mux_s11_h
    port map (
            O => \N__47005\,
            I => \N__47002\
        );

    \I__10243\ : Span12Mux_v
    port map (
            O => \N__47002\,
            I => \N__46999\
        );

    \I__10242\ : Odrv12
    port map (
            O => \N__46999\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__10241\ : InMux
    port map (
            O => \N__46996\,
            I => \N__46993\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__46993\,
            I => \N__46990\
        );

    \I__10239\ : Span4Mux_v
    port map (
            O => \N__46990\,
            I => \N__46986\
        );

    \I__10238\ : InMux
    port map (
            O => \N__46989\,
            I => \N__46983\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__46986\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__46983\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__10235\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46975\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__46975\,
            I => \N__46972\
        );

    \I__10233\ : Span4Mux_v
    port map (
            O => \N__46972\,
            I => \N__46968\
        );

    \I__10232\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46965\
        );

    \I__10231\ : Odrv4
    port map (
            O => \N__46968\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__46965\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__10229\ : InMux
    port map (
            O => \N__46960\,
            I => \N__46957\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__46957\,
            I => \N__46954\
        );

    \I__10227\ : Span4Mux_v
    port map (
            O => \N__46954\,
            I => \N__46950\
        );

    \I__10226\ : InMux
    port map (
            O => \N__46953\,
            I => \N__46947\
        );

    \I__10225\ : Odrv4
    port map (
            O => \N__46950\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__46947\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__10223\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46939\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__46939\,
            I => \N__46935\
        );

    \I__10221\ : InMux
    port map (
            O => \N__46938\,
            I => \N__46932\
        );

    \I__10220\ : Odrv12
    port map (
            O => \N__46935\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__46932\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10218\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46924\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__46924\,
            I => \N__46921\
        );

    \I__10216\ : Span4Mux_h
    port map (
            O => \N__46921\,
            I => \N__46917\
        );

    \I__10215\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46914\
        );

    \I__10214\ : Odrv4
    port map (
            O => \N__46917\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__46914\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__10212\ : CascadeMux
    port map (
            O => \N__46909\,
            I => \N__46905\
        );

    \I__10211\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46902\
        );

    \I__10210\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46899\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__46902\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__46899\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10207\ : InMux
    port map (
            O => \N__46894\,
            I => \N__46891\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__46891\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__10205\ : InMux
    port map (
            O => \N__46888\,
            I => \N__46885\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__46885\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__46882\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\
        );

    \I__10202\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46876\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__46876\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__10200\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46870\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__46870\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__46867\,
            I => \N__46864\
        );

    \I__10197\ : InMux
    port map (
            O => \N__46864\,
            I => \N__46858\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__46863\,
            I => \N__46855\
        );

    \I__10195\ : InMux
    port map (
            O => \N__46862\,
            I => \N__46852\
        );

    \I__10194\ : InMux
    port map (
            O => \N__46861\,
            I => \N__46849\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__46858\,
            I => \N__46846\
        );

    \I__10192\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46843\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__46852\,
            I => \N__46840\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__46849\,
            I => \N__46837\
        );

    \I__10189\ : Span4Mux_v
    port map (
            O => \N__46846\,
            I => \N__46832\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__46843\,
            I => \N__46832\
        );

    \I__10187\ : Span4Mux_h
    port map (
            O => \N__46840\,
            I => \N__46829\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__46837\,
            I => \N__46826\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__46832\,
            I => \N__46821\
        );

    \I__10184\ : Span4Mux_v
    port map (
            O => \N__46829\,
            I => \N__46821\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__46826\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10182\ : Odrv4
    port map (
            O => \N__46821\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__10181\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46813\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__46813\,
            I => \N__46810\
        );

    \I__10179\ : Span4Mux_h
    port map (
            O => \N__46810\,
            I => \N__46807\
        );

    \I__10178\ : Odrv4
    port map (
            O => \N__46807\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__10177\ : CascadeMux
    port map (
            O => \N__46804\,
            I => \N__46800\
        );

    \I__10176\ : InMux
    port map (
            O => \N__46803\,
            I => \N__46795\
        );

    \I__10175\ : InMux
    port map (
            O => \N__46800\,
            I => \N__46795\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__46795\,
            I => \N__46791\
        );

    \I__10173\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46788\
        );

    \I__10172\ : Span4Mux_h
    port map (
            O => \N__46791\,
            I => \N__46784\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__46788\,
            I => \N__46781\
        );

    \I__10170\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46778\
        );

    \I__10169\ : Odrv4
    port map (
            O => \N__46784\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__46781\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__46778\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__10166\ : InMux
    port map (
            O => \N__46771\,
            I => \N__46765\
        );

    \I__10165\ : InMux
    port map (
            O => \N__46770\,
            I => \N__46765\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__46765\,
            I => \N__46761\
        );

    \I__10163\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46758\
        );

    \I__10162\ : Odrv4
    port map (
            O => \N__46761\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__46758\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__10160\ : CascadeMux
    port map (
            O => \N__46753\,
            I => \N__46750\
        );

    \I__10159\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46747\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__46747\,
            I => \N__46744\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__46744\,
            I => \N__46741\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__46741\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__10155\ : InMux
    port map (
            O => \N__46738\,
            I => \N__46734\
        );

    \I__10154\ : InMux
    port map (
            O => \N__46737\,
            I => \N__46731\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__46734\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__46731\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__10151\ : InMux
    port map (
            O => \N__46726\,
            I => \N__46723\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__46723\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__10149\ : CascadeMux
    port map (
            O => \N__46720\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\
        );

    \I__10148\ : InMux
    port map (
            O => \N__46717\,
            I => \N__46714\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46711\
        );

    \I__10146\ : Span4Mux_v
    port map (
            O => \N__46711\,
            I => \N__46708\
        );

    \I__10145\ : Odrv4
    port map (
            O => \N__46708\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\
        );

    \I__10144\ : CascadeMux
    port map (
            O => \N__46705\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__10143\ : InMux
    port map (
            O => \N__46702\,
            I => \N__46699\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__46699\,
            I => \N__46695\
        );

    \I__10141\ : InMux
    port map (
            O => \N__46698\,
            I => \N__46692\
        );

    \I__10140\ : Span4Mux_v
    port map (
            O => \N__46695\,
            I => \N__46689\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__46692\,
            I => \N__46686\
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__46689\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__10137\ : Odrv4
    port map (
            O => \N__46686\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__10136\ : CascadeMux
    port map (
            O => \N__46681\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22_cascade_\
        );

    \I__10135\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46675\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__46675\,
            I => \N__46672\
        );

    \I__10133\ : Span4Mux_h
    port map (
            O => \N__46672\,
            I => \N__46669\
        );

    \I__10132\ : Odrv4
    port map (
            O => \N__46669\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__10131\ : CascadeMux
    port map (
            O => \N__46666\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__10130\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46660\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__46660\,
            I => \N__46656\
        );

    \I__10128\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46653\
        );

    \I__10127\ : Odrv4
    port map (
            O => \N__46656\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__46653\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__10125\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46644\
        );

    \I__10124\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46641\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46638\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46635\
        );

    \I__10121\ : Span4Mux_h
    port map (
            O => \N__46638\,
            I => \N__46632\
        );

    \I__10120\ : Odrv4
    port map (
            O => \N__46635\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10119\ : Odrv4
    port map (
            O => \N__46632\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10118\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46624\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__46624\,
            I => \N__46620\
        );

    \I__10116\ : InMux
    port map (
            O => \N__46623\,
            I => \N__46617\
        );

    \I__10115\ : Odrv4
    port map (
            O => \N__46620\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__46617\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__10113\ : InMux
    port map (
            O => \N__46612\,
            I => \N__46608\
        );

    \I__10112\ : InMux
    port map (
            O => \N__46611\,
            I => \N__46605\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__46608\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__46605\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__10109\ : InMux
    port map (
            O => \N__46600\,
            I => \N__46596\
        );

    \I__10108\ : CascadeMux
    port map (
            O => \N__46599\,
            I => \N__46593\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__46596\,
            I => \N__46590\
        );

    \I__10106\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46587\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__46590\,
            I => \N__46584\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__46587\,
            I => \N__46581\
        );

    \I__10103\ : Odrv4
    port map (
            O => \N__46584\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__10102\ : Odrv4
    port map (
            O => \N__46581\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__10101\ : InMux
    port map (
            O => \N__46576\,
            I => \N__46573\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__46573\,
            I => \N__46570\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__46570\,
            I => \N__46566\
        );

    \I__10098\ : InMux
    port map (
            O => \N__46569\,
            I => \N__46563\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__46566\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__46563\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10095\ : InMux
    port map (
            O => \N__46558\,
            I => \N__46554\
        );

    \I__10094\ : InMux
    port map (
            O => \N__46557\,
            I => \N__46551\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__46554\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__46551\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10091\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46543\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__46543\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__10089\ : CascadeMux
    port map (
            O => \N__46540\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\
        );

    \I__10088\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46534\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__46534\,
            I => \N__46531\
        );

    \I__10086\ : Span4Mux_v
    port map (
            O => \N__46531\,
            I => \N__46528\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__46528\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\
        );

    \I__10084\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46509\
        );

    \I__10083\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46509\
        );

    \I__10082\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46509\
        );

    \I__10081\ : InMux
    port map (
            O => \N__46522\,
            I => \N__46509\
        );

    \I__10080\ : InMux
    port map (
            O => \N__46521\,
            I => \N__46490\
        );

    \I__10079\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46490\
        );

    \I__10078\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46490\
        );

    \I__10077\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46490\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__46509\,
            I => \N__46487\
        );

    \I__10075\ : InMux
    port map (
            O => \N__46508\,
            I => \N__46478\
        );

    \I__10074\ : InMux
    port map (
            O => \N__46507\,
            I => \N__46478\
        );

    \I__10073\ : InMux
    port map (
            O => \N__46506\,
            I => \N__46478\
        );

    \I__10072\ : InMux
    port map (
            O => \N__46505\,
            I => \N__46478\
        );

    \I__10071\ : InMux
    port map (
            O => \N__46504\,
            I => \N__46469\
        );

    \I__10070\ : InMux
    port map (
            O => \N__46503\,
            I => \N__46469\
        );

    \I__10069\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46469\
        );

    \I__10068\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46469\
        );

    \I__10067\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46452\
        );

    \I__10066\ : InMux
    port map (
            O => \N__46499\,
            I => \N__46452\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__46490\,
            I => \N__46443\
        );

    \I__10064\ : Span4Mux_h
    port map (
            O => \N__46487\,
            I => \N__46443\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__46478\,
            I => \N__46443\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__46469\,
            I => \N__46443\
        );

    \I__10061\ : InMux
    port map (
            O => \N__46468\,
            I => \N__46434\
        );

    \I__10060\ : InMux
    port map (
            O => \N__46467\,
            I => \N__46434\
        );

    \I__10059\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46434\
        );

    \I__10058\ : InMux
    port map (
            O => \N__46465\,
            I => \N__46434\
        );

    \I__10057\ : InMux
    port map (
            O => \N__46464\,
            I => \N__46425\
        );

    \I__10056\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46425\
        );

    \I__10055\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46425\
        );

    \I__10054\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46425\
        );

    \I__10053\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46416\
        );

    \I__10052\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46416\
        );

    \I__10051\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46416\
        );

    \I__10050\ : InMux
    port map (
            O => \N__46457\,
            I => \N__46416\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__46452\,
            I => \N__46413\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__46443\,
            I => \N__46410\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__46434\,
            I => \N__46403\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__46425\,
            I => \N__46403\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__46416\,
            I => \N__46403\
        );

    \I__10044\ : Odrv4
    port map (
            O => \N__46413\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__10043\ : Odrv4
    port map (
            O => \N__46410\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__10042\ : Odrv12
    port map (
            O => \N__46403\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__10041\ : CascadeMux
    port map (
            O => \N__46396\,
            I => \N__46393\
        );

    \I__10040\ : InMux
    port map (
            O => \N__46393\,
            I => \N__46389\
        );

    \I__10039\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46386\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__46389\,
            I => \N__46380\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__46386\,
            I => \N__46380\
        );

    \I__10036\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46377\
        );

    \I__10035\ : Span4Mux_h
    port map (
            O => \N__46380\,
            I => \N__46374\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__46377\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__46374\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10032\ : InMux
    port map (
            O => \N__46369\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__10031\ : CascadeMux
    port map (
            O => \N__46366\,
            I => \N__46363\
        );

    \I__10030\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46359\
        );

    \I__10029\ : InMux
    port map (
            O => \N__46362\,
            I => \N__46356\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46350\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__46356\,
            I => \N__46350\
        );

    \I__10026\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46347\
        );

    \I__10025\ : Span4Mux_h
    port map (
            O => \N__46350\,
            I => \N__46344\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__46347\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10023\ : Odrv4
    port map (
            O => \N__46344\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10022\ : InMux
    port map (
            O => \N__46339\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__10021\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46333\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__46333\,
            I => \N__46329\
        );

    \I__10019\ : InMux
    port map (
            O => \N__46332\,
            I => \N__46326\
        );

    \I__10018\ : Span4Mux_h
    port map (
            O => \N__46329\,
            I => \N__46323\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__46326\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10016\ : Odrv4
    port map (
            O => \N__46323\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10015\ : InMux
    port map (
            O => \N__46318\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__10014\ : InMux
    port map (
            O => \N__46315\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__10013\ : InMux
    port map (
            O => \N__46312\,
            I => \N__46308\
        );

    \I__10012\ : InMux
    port map (
            O => \N__46311\,
            I => \N__46305\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__46308\,
            I => \N__46302\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__46305\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10009\ : Odrv4
    port map (
            O => \N__46302\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10008\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46294\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46291\
        );

    \I__10006\ : Span4Mux_v
    port map (
            O => \N__46291\,
            I => \N__46287\
        );

    \I__10005\ : InMux
    port map (
            O => \N__46290\,
            I => \N__46284\
        );

    \I__10004\ : Odrv4
    port map (
            O => \N__46287\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__46284\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10002\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46276\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__46276\,
            I => \N__46272\
        );

    \I__10000\ : InMux
    port map (
            O => \N__46275\,
            I => \N__46269\
        );

    \I__9999\ : Odrv4
    port map (
            O => \N__46272\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__46269\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__9997\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46260\
        );

    \I__9996\ : CascadeMux
    port map (
            O => \N__46263\,
            I => \N__46257\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__46260\,
            I => \N__46254\
        );

    \I__9994\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46251\
        );

    \I__9993\ : Odrv4
    port map (
            O => \N__46254\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__46251\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__9991\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46243\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__46243\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__9989\ : CascadeMux
    port map (
            O => \N__46240\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__9988\ : InMux
    port map (
            O => \N__46237\,
            I => \N__46234\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__46234\,
            I => \N__46231\
        );

    \I__9986\ : Odrv12
    port map (
            O => \N__46231\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\
        );

    \I__9985\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46225\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__46225\,
            I => \N__46221\
        );

    \I__9983\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46218\
        );

    \I__9982\ : Odrv4
    port map (
            O => \N__46221\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__46218\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9980\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46210\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__46210\,
            I => \N__46206\
        );

    \I__9978\ : InMux
    port map (
            O => \N__46209\,
            I => \N__46203\
        );

    \I__9977\ : Odrv4
    port map (
            O => \N__46206\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__46203\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__9975\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46194\
        );

    \I__9974\ : CascadeMux
    port map (
            O => \N__46197\,
            I => \N__46191\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__46194\,
            I => \N__46188\
        );

    \I__9972\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46185\
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__46188\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__46185\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9969\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46177\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__46177\,
            I => \N__46173\
        );

    \I__9967\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46170\
        );

    \I__9966\ : Odrv4
    port map (
            O => \N__46173\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__46170\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__9964\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46159\
        );

    \I__9963\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46159\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__46159\,
            I => \N__46155\
        );

    \I__9961\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46152\
        );

    \I__9960\ : Span4Mux_h
    port map (
            O => \N__46155\,
            I => \N__46149\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__46152\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__46149\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9957\ : InMux
    port map (
            O => \N__46144\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__9956\ : InMux
    port map (
            O => \N__46141\,
            I => \N__46134\
        );

    \I__9955\ : InMux
    port map (
            O => \N__46140\,
            I => \N__46134\
        );

    \I__9954\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46131\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__46134\,
            I => \N__46128\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__46131\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9951\ : Odrv4
    port map (
            O => \N__46128\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9950\ : InMux
    port map (
            O => \N__46123\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__9949\ : CascadeMux
    port map (
            O => \N__46120\,
            I => \N__46116\
        );

    \I__9948\ : CascadeMux
    port map (
            O => \N__46119\,
            I => \N__46113\
        );

    \I__9947\ : InMux
    port map (
            O => \N__46116\,
            I => \N__46107\
        );

    \I__9946\ : InMux
    port map (
            O => \N__46113\,
            I => \N__46107\
        );

    \I__9945\ : InMux
    port map (
            O => \N__46112\,
            I => \N__46104\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__46107\,
            I => \N__46101\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__46104\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9942\ : Odrv4
    port map (
            O => \N__46101\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9941\ : InMux
    port map (
            O => \N__46096\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__46093\,
            I => \N__46090\
        );

    \I__9939\ : InMux
    port map (
            O => \N__46090\,
            I => \N__46086\
        );

    \I__9938\ : InMux
    port map (
            O => \N__46089\,
            I => \N__46082\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__46079\
        );

    \I__9936\ : InMux
    port map (
            O => \N__46085\,
            I => \N__46076\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__46082\,
            I => \N__46071\
        );

    \I__9934\ : Span4Mux_h
    port map (
            O => \N__46079\,
            I => \N__46071\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__46076\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9932\ : Odrv4
    port map (
            O => \N__46071\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9931\ : InMux
    port map (
            O => \N__46066\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__9930\ : InMux
    port map (
            O => \N__46063\,
            I => \N__46056\
        );

    \I__9929\ : InMux
    port map (
            O => \N__46062\,
            I => \N__46056\
        );

    \I__9928\ : InMux
    port map (
            O => \N__46061\,
            I => \N__46053\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__46056\,
            I => \N__46050\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__46053\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__46050\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9924\ : InMux
    port map (
            O => \N__46045\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__9923\ : CascadeMux
    port map (
            O => \N__46042\,
            I => \N__46038\
        );

    \I__9922\ : CascadeMux
    port map (
            O => \N__46041\,
            I => \N__46035\
        );

    \I__9921\ : InMux
    port map (
            O => \N__46038\,
            I => \N__46029\
        );

    \I__9920\ : InMux
    port map (
            O => \N__46035\,
            I => \N__46029\
        );

    \I__9919\ : InMux
    port map (
            O => \N__46034\,
            I => \N__46026\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__46029\,
            I => \N__46023\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__46026\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9916\ : Odrv4
    port map (
            O => \N__46023\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9915\ : InMux
    port map (
            O => \N__46018\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__9914\ : CascadeMux
    port map (
            O => \N__46015\,
            I => \N__46012\
        );

    \I__9913\ : InMux
    port map (
            O => \N__46012\,
            I => \N__46007\
        );

    \I__9912\ : CascadeMux
    port map (
            O => \N__46011\,
            I => \N__46004\
        );

    \I__9911\ : InMux
    port map (
            O => \N__46010\,
            I => \N__46001\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__46007\,
            I => \N__45998\
        );

    \I__9909\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45995\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__46001\,
            I => \N__45990\
        );

    \I__9907\ : Span4Mux_v
    port map (
            O => \N__45998\,
            I => \N__45990\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__45995\,
            I => \N__45987\
        );

    \I__9905\ : Odrv4
    port map (
            O => \N__45990\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9904\ : Odrv4
    port map (
            O => \N__45987\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9903\ : InMux
    port map (
            O => \N__45982\,
            I => \bfn_18_10_0_\
        );

    \I__9902\ : CascadeMux
    port map (
            O => \N__45979\,
            I => \N__45976\
        );

    \I__9901\ : InMux
    port map (
            O => \N__45976\,
            I => \N__45973\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__45973\,
            I => \N__45968\
        );

    \I__9899\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45965\
        );

    \I__9898\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45962\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__45968\,
            I => \N__45959\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45956\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__45962\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9894\ : Odrv4
    port map (
            O => \N__45959\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9893\ : Odrv4
    port map (
            O => \N__45956\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9892\ : InMux
    port map (
            O => \N__45949\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__9891\ : CascadeMux
    port map (
            O => \N__45946\,
            I => \N__45943\
        );

    \I__9890\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45938\
        );

    \I__9889\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45935\
        );

    \I__9888\ : InMux
    port map (
            O => \N__45941\,
            I => \N__45932\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__45938\,
            I => \N__45929\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__45935\,
            I => \N__45926\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__45932\,
            I => \N__45921\
        );

    \I__9884\ : Span4Mux_v
    port map (
            O => \N__45929\,
            I => \N__45921\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__45926\,
            I => \N__45918\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__45921\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__45918\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9880\ : InMux
    port map (
            O => \N__45913\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__9879\ : CascadeMux
    port map (
            O => \N__45910\,
            I => \N__45906\
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__45909\,
            I => \N__45903\
        );

    \I__9877\ : InMux
    port map (
            O => \N__45906\,
            I => \N__45897\
        );

    \I__9876\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45897\
        );

    \I__9875\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45894\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45891\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__45894\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9872\ : Odrv4
    port map (
            O => \N__45891\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9871\ : InMux
    port map (
            O => \N__45886\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__9870\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45877\
        );

    \I__9869\ : InMux
    port map (
            O => \N__45882\,
            I => \N__45877\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__45877\,
            I => \N__45873\
        );

    \I__9867\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45870\
        );

    \I__9866\ : Span4Mux_h
    port map (
            O => \N__45873\,
            I => \N__45867\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__45870\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9864\ : Odrv4
    port map (
            O => \N__45867\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9863\ : InMux
    port map (
            O => \N__45862\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__9862\ : CascadeMux
    port map (
            O => \N__45859\,
            I => \N__45856\
        );

    \I__9861\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45852\
        );

    \I__9860\ : InMux
    port map (
            O => \N__45855\,
            I => \N__45849\
        );

    \I__9859\ : LocalMux
    port map (
            O => \N__45852\,
            I => \N__45843\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__45849\,
            I => \N__45843\
        );

    \I__9857\ : InMux
    port map (
            O => \N__45848\,
            I => \N__45840\
        );

    \I__9856\ : Span4Mux_h
    port map (
            O => \N__45843\,
            I => \N__45837\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__45840\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__45837\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9853\ : InMux
    port map (
            O => \N__45832\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__45829\,
            I => \N__45826\
        );

    \I__9851\ : InMux
    port map (
            O => \N__45826\,
            I => \N__45822\
        );

    \I__9850\ : InMux
    port map (
            O => \N__45825\,
            I => \N__45818\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__45822\,
            I => \N__45815\
        );

    \I__9848\ : InMux
    port map (
            O => \N__45821\,
            I => \N__45812\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__45818\,
            I => \N__45807\
        );

    \I__9846\ : Span4Mux_h
    port map (
            O => \N__45815\,
            I => \N__45807\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__45812\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9844\ : Odrv4
    port map (
            O => \N__45807\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9843\ : InMux
    port map (
            O => \N__45802\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__9842\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45792\
        );

    \I__9841\ : InMux
    port map (
            O => \N__45798\,
            I => \N__45792\
        );

    \I__9840\ : InMux
    port map (
            O => \N__45797\,
            I => \N__45789\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__45792\,
            I => \N__45786\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__45789\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__45786\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9836\ : InMux
    port map (
            O => \N__45781\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__9835\ : CascadeMux
    port map (
            O => \N__45778\,
            I => \N__45774\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__45777\,
            I => \N__45771\
        );

    \I__9833\ : InMux
    port map (
            O => \N__45774\,
            I => \N__45765\
        );

    \I__9832\ : InMux
    port map (
            O => \N__45771\,
            I => \N__45765\
        );

    \I__9831\ : InMux
    port map (
            O => \N__45770\,
            I => \N__45762\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45759\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__45762\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9828\ : Odrv4
    port map (
            O => \N__45759\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9827\ : InMux
    port map (
            O => \N__45754\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__45751\,
            I => \N__45748\
        );

    \I__9825\ : InMux
    port map (
            O => \N__45748\,
            I => \N__45744\
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__45747\,
            I => \N__45741\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__45744\,
            I => \N__45737\
        );

    \I__9822\ : InMux
    port map (
            O => \N__45741\,
            I => \N__45734\
        );

    \I__9821\ : InMux
    port map (
            O => \N__45740\,
            I => \N__45731\
        );

    \I__9820\ : Span4Mux_v
    port map (
            O => \N__45737\,
            I => \N__45726\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__45734\,
            I => \N__45726\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__45731\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9817\ : Odrv4
    port map (
            O => \N__45726\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9816\ : InMux
    port map (
            O => \N__45721\,
            I => \bfn_18_9_0_\
        );

    \I__9815\ : CascadeMux
    port map (
            O => \N__45718\,
            I => \N__45715\
        );

    \I__9814\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45712\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__45712\,
            I => \N__45707\
        );

    \I__9812\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45704\
        );

    \I__9811\ : InMux
    port map (
            O => \N__45710\,
            I => \N__45701\
        );

    \I__9810\ : Span4Mux_v
    port map (
            O => \N__45707\,
            I => \N__45698\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__45704\,
            I => \N__45695\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__45701\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9807\ : Odrv4
    port map (
            O => \N__45698\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__45695\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9805\ : InMux
    port map (
            O => \N__45688\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__9804\ : InMux
    port map (
            O => \N__45685\,
            I => \N__45681\
        );

    \I__9803\ : CascadeMux
    port map (
            O => \N__45684\,
            I => \N__45678\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__45681\,
            I => \N__45674\
        );

    \I__9801\ : InMux
    port map (
            O => \N__45678\,
            I => \N__45671\
        );

    \I__9800\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45668\
        );

    \I__9799\ : Span4Mux_h
    port map (
            O => \N__45674\,
            I => \N__45663\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__45671\,
            I => \N__45663\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__45668\,
            I => \N__45658\
        );

    \I__9796\ : Span4Mux_v
    port map (
            O => \N__45663\,
            I => \N__45658\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__45658\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9794\ : InMux
    port map (
            O => \N__45655\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__9793\ : CascadeMux
    port map (
            O => \N__45652\,
            I => \N__45648\
        );

    \I__9792\ : CascadeMux
    port map (
            O => \N__45651\,
            I => \N__45645\
        );

    \I__9791\ : InMux
    port map (
            O => \N__45648\,
            I => \N__45639\
        );

    \I__9790\ : InMux
    port map (
            O => \N__45645\,
            I => \N__45639\
        );

    \I__9789\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45636\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__45639\,
            I => \N__45633\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__45636\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9786\ : Odrv4
    port map (
            O => \N__45633\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9785\ : InMux
    port map (
            O => \N__45628\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__9784\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45618\
        );

    \I__9783\ : InMux
    port map (
            O => \N__45624\,
            I => \N__45618\
        );

    \I__9782\ : InMux
    port map (
            O => \N__45623\,
            I => \N__45615\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__45618\,
            I => \N__45612\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__45615\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9779\ : Odrv4
    port map (
            O => \N__45612\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9778\ : InMux
    port map (
            O => \N__45607\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__9777\ : CascadeMux
    port map (
            O => \N__45604\,
            I => \N__45600\
        );

    \I__9776\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45597\
        );

    \I__9775\ : InMux
    port map (
            O => \N__45600\,
            I => \N__45593\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__45597\,
            I => \N__45590\
        );

    \I__9773\ : InMux
    port map (
            O => \N__45596\,
            I => \N__45587\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__45593\,
            I => \N__45582\
        );

    \I__9771\ : Span4Mux_h
    port map (
            O => \N__45590\,
            I => \N__45582\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__45587\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9769\ : Odrv4
    port map (
            O => \N__45582\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9768\ : InMux
    port map (
            O => \N__45577\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__9767\ : CascadeMux
    port map (
            O => \N__45574\,
            I => \N__45570\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__45573\,
            I => \N__45567\
        );

    \I__9765\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45562\
        );

    \I__9764\ : InMux
    port map (
            O => \N__45567\,
            I => \N__45562\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__45562\,
            I => \N__45558\
        );

    \I__9762\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45555\
        );

    \I__9761\ : Span4Mux_h
    port map (
            O => \N__45558\,
            I => \N__45552\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__45555\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9759\ : Odrv4
    port map (
            O => \N__45552\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9758\ : InMux
    port map (
            O => \N__45547\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45537\
        );

    \I__9756\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45537\
        );

    \I__9755\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45534\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__45537\,
            I => \N__45531\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__45534\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9752\ : Odrv4
    port map (
            O => \N__45531\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9751\ : InMux
    port map (
            O => \N__45526\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__9750\ : CascadeMux
    port map (
            O => \N__45523\,
            I => \N__45520\
        );

    \I__9749\ : InMux
    port map (
            O => \N__45520\,
            I => \N__45516\
        );

    \I__9748\ : InMux
    port map (
            O => \N__45519\,
            I => \N__45513\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__45516\,
            I => \N__45507\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__45513\,
            I => \N__45507\
        );

    \I__9745\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45504\
        );

    \I__9744\ : Span4Mux_h
    port map (
            O => \N__45507\,
            I => \N__45501\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__45504\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9742\ : Odrv4
    port map (
            O => \N__45501\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9741\ : InMux
    port map (
            O => \N__45496\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__9740\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45489\
        );

    \I__9739\ : CascadeMux
    port map (
            O => \N__45492\,
            I => \N__45486\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__45489\,
            I => \N__45482\
        );

    \I__9737\ : InMux
    port map (
            O => \N__45486\,
            I => \N__45479\
        );

    \I__9736\ : InMux
    port map (
            O => \N__45485\,
            I => \N__45476\
        );

    \I__9735\ : Span4Mux_v
    port map (
            O => \N__45482\,
            I => \N__45471\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__45479\,
            I => \N__45471\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__45476\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__45471\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9731\ : InMux
    port map (
            O => \N__45466\,
            I => \bfn_18_8_0_\
        );

    \I__9730\ : CascadeMux
    port map (
            O => \N__45463\,
            I => \N__45460\
        );

    \I__9729\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45457\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__45457\,
            I => \N__45454\
        );

    \I__9727\ : Odrv4
    port map (
            O => \N__45454\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__9726\ : InMux
    port map (
            O => \N__45451\,
            I => \N__45448\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__45448\,
            I => \N__45445\
        );

    \I__9724\ : Span4Mux_h
    port map (
            O => \N__45445\,
            I => \N__45442\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__45442\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__9722\ : InMux
    port map (
            O => \N__45439\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__9721\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45433\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__45433\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__9719\ : InMux
    port map (
            O => \N__45430\,
            I => \N__45427\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__45427\,
            I => \N__45424\
        );

    \I__9717\ : Odrv12
    port map (
            O => \N__45424\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__9716\ : InMux
    port map (
            O => \N__45421\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__9715\ : CascadeMux
    port map (
            O => \N__45418\,
            I => \N__45415\
        );

    \I__9714\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45412\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__45412\,
            I => \N__45409\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__45409\,
            I => \N__45406\
        );

    \I__9711\ : Span4Mux_v
    port map (
            O => \N__45406\,
            I => \N__45403\
        );

    \I__9710\ : Span4Mux_v
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__9709\ : Odrv4
    port map (
            O => \N__45400\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__9708\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45394\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__45394\,
            I => \N__45391\
        );

    \I__9706\ : Odrv4
    port map (
            O => \N__45391\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__9705\ : InMux
    port map (
            O => \N__45388\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__9704\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45382\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__45382\,
            I => \N__45379\
        );

    \I__9702\ : Span4Mux_v
    port map (
            O => \N__45379\,
            I => \N__45376\
        );

    \I__9701\ : Span4Mux_v
    port map (
            O => \N__45376\,
            I => \N__45373\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__45373\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__9699\ : InMux
    port map (
            O => \N__45370\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__9698\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45364\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45361\
        );

    \I__9696\ : Span4Mux_h
    port map (
            O => \N__45361\,
            I => \N__45358\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__45358\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__9694\ : InMux
    port map (
            O => \N__45355\,
            I => \N__45352\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__45352\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__45349\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\
        );

    \I__9691\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45343\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__45343\,
            I => \N__45340\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__45340\,
            I => \N__45337\
        );

    \I__9688\ : Span4Mux_v
    port map (
            O => \N__45337\,
            I => \N__45334\
        );

    \I__9687\ : Odrv4
    port map (
            O => \N__45334\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\
        );

    \I__9686\ : InMux
    port map (
            O => \N__45331\,
            I => \N__45327\
        );

    \I__9685\ : InMux
    port map (
            O => \N__45330\,
            I => \N__45324\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__45327\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__45324\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__9682\ : InMux
    port map (
            O => \N__45319\,
            I => \N__45316\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__45316\,
            I => \N__45312\
        );

    \I__9680\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45309\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__45312\,
            I => \N__45304\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__45309\,
            I => \N__45304\
        );

    \I__9677\ : Span4Mux_v
    port map (
            O => \N__45304\,
            I => \N__45300\
        );

    \I__9676\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45297\
        );

    \I__9675\ : Odrv4
    port map (
            O => \N__45300\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__45297\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9673\ : InMux
    port map (
            O => \N__45292\,
            I => \bfn_18_7_0_\
        );

    \I__9672\ : CascadeMux
    port map (
            O => \N__45289\,
            I => \N__45286\
        );

    \I__9671\ : InMux
    port map (
            O => \N__45286\,
            I => \N__45283\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__45283\,
            I => \N__45280\
        );

    \I__9669\ : Odrv12
    port map (
            O => \N__45280\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__9668\ : InMux
    port map (
            O => \N__45277\,
            I => \N__45274\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__45274\,
            I => \N__45271\
        );

    \I__9666\ : Span4Mux_v
    port map (
            O => \N__45271\,
            I => \N__45268\
        );

    \I__9665\ : Sp12to4
    port map (
            O => \N__45268\,
            I => \N__45265\
        );

    \I__9664\ : Odrv12
    port map (
            O => \N__45265\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__9663\ : InMux
    port map (
            O => \N__45262\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__9662\ : InMux
    port map (
            O => \N__45259\,
            I => \N__45256\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__45256\,
            I => \N__45253\
        );

    \I__9660\ : Odrv12
    port map (
            O => \N__45253\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__9659\ : InMux
    port map (
            O => \N__45250\,
            I => \N__45247\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45244\
        );

    \I__9657\ : Span4Mux_v
    port map (
            O => \N__45244\,
            I => \N__45241\
        );

    \I__9656\ : Sp12to4
    port map (
            O => \N__45241\,
            I => \N__45238\
        );

    \I__9655\ : Odrv12
    port map (
            O => \N__45238\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__9654\ : InMux
    port map (
            O => \N__45235\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__45232\,
            I => \N__45229\
        );

    \I__9652\ : InMux
    port map (
            O => \N__45229\,
            I => \N__45226\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__45226\,
            I => \N__45223\
        );

    \I__9650\ : Span4Mux_h
    port map (
            O => \N__45223\,
            I => \N__45220\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__45220\,
            I => \N__45217\
        );

    \I__9648\ : Odrv4
    port map (
            O => \N__45217\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__9647\ : InMux
    port map (
            O => \N__45214\,
            I => \N__45211\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__45211\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__9645\ : InMux
    port map (
            O => \N__45208\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__9644\ : InMux
    port map (
            O => \N__45205\,
            I => \N__45202\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__45202\,
            I => \N__45199\
        );

    \I__9642\ : Odrv12
    port map (
            O => \N__45199\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__9641\ : InMux
    port map (
            O => \N__45196\,
            I => \N__45193\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__45193\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__9639\ : InMux
    port map (
            O => \N__45190\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__9638\ : CascadeMux
    port map (
            O => \N__45187\,
            I => \N__45184\
        );

    \I__9637\ : InMux
    port map (
            O => \N__45184\,
            I => \N__45181\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__45181\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__9635\ : InMux
    port map (
            O => \N__45178\,
            I => \N__45175\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__45175\,
            I => \N__45172\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__45172\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__9632\ : InMux
    port map (
            O => \N__45169\,
            I => \bfn_17_21_0_\
        );

    \I__9631\ : InMux
    port map (
            O => \N__45166\,
            I => \N__45163\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__45163\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__9629\ : InMux
    port map (
            O => \N__45160\,
            I => \N__45157\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__45157\,
            I => \N__45154\
        );

    \I__9627\ : Odrv4
    port map (
            O => \N__45154\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__9626\ : InMux
    port map (
            O => \N__45151\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__9625\ : CascadeMux
    port map (
            O => \N__45148\,
            I => \N__45145\
        );

    \I__9624\ : InMux
    port map (
            O => \N__45145\,
            I => \N__45142\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__45142\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__9622\ : InMux
    port map (
            O => \N__45139\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__9621\ : InMux
    port map (
            O => \N__45136\,
            I => \N__45133\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__45133\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__9619\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45127\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__45127\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__9617\ : InMux
    port map (
            O => \N__45124\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__45121\,
            I => \N__45118\
        );

    \I__9615\ : InMux
    port map (
            O => \N__45118\,
            I => \N__45115\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__45115\,
            I => \N__45112\
        );

    \I__9613\ : Odrv12
    port map (
            O => \N__45112\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__9612\ : InMux
    port map (
            O => \N__45109\,
            I => \N__45106\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__45106\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__9610\ : InMux
    port map (
            O => \N__45103\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__9609\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45097\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__45097\,
            I => \N__45094\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__45094\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__9606\ : InMux
    port map (
            O => \N__45091\,
            I => \N__45088\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__45088\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__9604\ : InMux
    port map (
            O => \N__45085\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__45082\,
            I => \N__45079\
        );

    \I__9602\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45076\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__45076\,
            I => \N__45073\
        );

    \I__9600\ : Odrv12
    port map (
            O => \N__45073\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__9599\ : InMux
    port map (
            O => \N__45070\,
            I => \N__45067\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__45067\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__9597\ : InMux
    port map (
            O => \N__45064\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__9596\ : InMux
    port map (
            O => \N__45061\,
            I => \N__45058\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__45058\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__9594\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45052\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__45052\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__9592\ : InMux
    port map (
            O => \N__45049\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__9591\ : CascadeMux
    port map (
            O => \N__45046\,
            I => \N__45043\
        );

    \I__9590\ : InMux
    port map (
            O => \N__45043\,
            I => \N__45040\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__45040\,
            I => \N__45037\
        );

    \I__9588\ : Odrv12
    port map (
            O => \N__45037\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__9587\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45031\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__45031\,
            I => \N__45028\
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__45028\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__9584\ : InMux
    port map (
            O => \N__45025\,
            I => \bfn_17_20_0_\
        );

    \I__9583\ : InMux
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__45019\,
            I => \N__45016\
        );

    \I__9581\ : Span4Mux_v
    port map (
            O => \N__45016\,
            I => \N__45013\
        );

    \I__9580\ : Odrv4
    port map (
            O => \N__45013\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__9579\ : InMux
    port map (
            O => \N__45010\,
            I => \N__45007\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__45007\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__9577\ : InMux
    port map (
            O => \N__45004\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__9576\ : CascadeMux
    port map (
            O => \N__45001\,
            I => \N__44998\
        );

    \I__9575\ : InMux
    port map (
            O => \N__44998\,
            I => \N__44995\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__44995\,
            I => \N__44992\
        );

    \I__9573\ : Span12Mux_s9_h
    port map (
            O => \N__44992\,
            I => \N__44989\
        );

    \I__9572\ : Odrv12
    port map (
            O => \N__44989\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__9571\ : InMux
    port map (
            O => \N__44986\,
            I => \N__44983\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__44983\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__9569\ : InMux
    port map (
            O => \N__44980\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__9568\ : InMux
    port map (
            O => \N__44977\,
            I => \N__44974\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__44974\,
            I => \N__44971\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__44971\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__9565\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44965\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__44965\,
            I => \N__44962\
        );

    \I__9563\ : Span4Mux_h
    port map (
            O => \N__44962\,
            I => \N__44959\
        );

    \I__9562\ : Odrv4
    port map (
            O => \N__44959\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__9561\ : InMux
    port map (
            O => \N__44956\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__9560\ : CascadeMux
    port map (
            O => \N__44953\,
            I => \N__44950\
        );

    \I__9559\ : InMux
    port map (
            O => \N__44950\,
            I => \N__44947\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__44947\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__9557\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44941\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__44941\,
            I => \N__44938\
        );

    \I__9555\ : Span4Mux_h
    port map (
            O => \N__44938\,
            I => \N__44935\
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__44935\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__9553\ : InMux
    port map (
            O => \N__44932\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__9552\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44926\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__44926\,
            I => \N__44923\
        );

    \I__9550\ : Span4Mux_v
    port map (
            O => \N__44923\,
            I => \N__44920\
        );

    \I__9549\ : Odrv4
    port map (
            O => \N__44920\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__9548\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44914\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__44914\,
            I => \N__44911\
        );

    \I__9546\ : Span4Mux_v
    port map (
            O => \N__44911\,
            I => \N__44908\
        );

    \I__9545\ : Odrv4
    port map (
            O => \N__44908\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__9544\ : InMux
    port map (
            O => \N__44905\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__9543\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44899\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44896\
        );

    \I__9541\ : Span4Mux_v
    port map (
            O => \N__44896\,
            I => \N__44893\
        );

    \I__9540\ : Odrv4
    port map (
            O => \N__44893\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__9539\ : InMux
    port map (
            O => \N__44890\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__9538\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44884\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__44884\,
            I => \N__44881\
        );

    \I__9536\ : Span4Mux_h
    port map (
            O => \N__44881\,
            I => \N__44878\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__44878\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__9534\ : InMux
    port map (
            O => \N__44875\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__9533\ : CascadeMux
    port map (
            O => \N__44872\,
            I => \N__44869\
        );

    \I__9532\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44866\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__44866\,
            I => \N__44863\
        );

    \I__9530\ : Span4Mux_v
    port map (
            O => \N__44863\,
            I => \N__44860\
        );

    \I__9529\ : Odrv4
    port map (
            O => \N__44860\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__9528\ : InMux
    port map (
            O => \N__44857\,
            I => \N__44854\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__44854\,
            I => \N__44851\
        );

    \I__9526\ : Span4Mux_v
    port map (
            O => \N__44851\,
            I => \N__44848\
        );

    \I__9525\ : Odrv4
    port map (
            O => \N__44848\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__9524\ : InMux
    port map (
            O => \N__44845\,
            I => \bfn_17_19_0_\
        );

    \I__9523\ : InMux
    port map (
            O => \N__44842\,
            I => \N__44839\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__44839\,
            I => \N__44836\
        );

    \I__9521\ : Odrv12
    port map (
            O => \N__44836\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__9520\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44830\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__44830\,
            I => \N__44827\
        );

    \I__9518\ : Span4Mux_h
    port map (
            O => \N__44827\,
            I => \N__44824\
        );

    \I__9517\ : Odrv4
    port map (
            O => \N__44824\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__9516\ : InMux
    port map (
            O => \N__44821\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__44818\,
            I => \N__44815\
        );

    \I__9514\ : InMux
    port map (
            O => \N__44815\,
            I => \N__44812\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__44812\,
            I => \N__44809\
        );

    \I__9512\ : Span4Mux_v
    port map (
            O => \N__44809\,
            I => \N__44806\
        );

    \I__9511\ : Odrv4
    port map (
            O => \N__44806\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__9510\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44800\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__44800\,
            I => \N__44797\
        );

    \I__9508\ : Span4Mux_v
    port map (
            O => \N__44797\,
            I => \N__44794\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__44794\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__9506\ : InMux
    port map (
            O => \N__44791\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__9505\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44785\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__44785\,
            I => \N__44782\
        );

    \I__9503\ : Odrv12
    port map (
            O => \N__44782\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__9502\ : InMux
    port map (
            O => \N__44779\,
            I => \N__44776\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__44776\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__9500\ : InMux
    port map (
            O => \N__44773\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__9499\ : CascadeMux
    port map (
            O => \N__44770\,
            I => \N__44767\
        );

    \I__9498\ : InMux
    port map (
            O => \N__44767\,
            I => \N__44762\
        );

    \I__9497\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44756\
        );

    \I__9496\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44756\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__44762\,
            I => \N__44753\
        );

    \I__9494\ : InMux
    port map (
            O => \N__44761\,
            I => \N__44750\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__44756\,
            I => \N__44747\
        );

    \I__9492\ : Span4Mux_v
    port map (
            O => \N__44753\,
            I => \N__44744\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__44750\,
            I => \N__44741\
        );

    \I__9490\ : Span4Mux_h
    port map (
            O => \N__44747\,
            I => \N__44738\
        );

    \I__9489\ : Odrv4
    port map (
            O => \N__44744\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9488\ : Odrv12
    port map (
            O => \N__44741\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9487\ : Odrv4
    port map (
            O => \N__44738\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9486\ : InMux
    port map (
            O => \N__44731\,
            I => \N__44727\
        );

    \I__9485\ : CascadeMux
    port map (
            O => \N__44730\,
            I => \N__44724\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__44727\,
            I => \N__44720\
        );

    \I__9483\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44717\
        );

    \I__9482\ : InMux
    port map (
            O => \N__44723\,
            I => \N__44714\
        );

    \I__9481\ : Odrv12
    port map (
            O => \N__44720\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__44717\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__44714\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9478\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44700\
        );

    \I__9477\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44700\
        );

    \I__9476\ : CascadeMux
    port map (
            O => \N__44705\,
            I => \N__44697\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__44700\,
            I => \N__44694\
        );

    \I__9474\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44691\
        );

    \I__9473\ : Span4Mux_h
    port map (
            O => \N__44694\,
            I => \N__44688\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__44691\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9471\ : Odrv4
    port map (
            O => \N__44688\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9470\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44677\
        );

    \I__9469\ : InMux
    port map (
            O => \N__44682\,
            I => \N__44677\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__44677\,
            I => \N__44673\
        );

    \I__9467\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44670\
        );

    \I__9466\ : Span4Mux_h
    port map (
            O => \N__44673\,
            I => \N__44664\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__44670\,
            I => \N__44664\
        );

    \I__9464\ : InMux
    port map (
            O => \N__44669\,
            I => \N__44661\
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__44664\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__44661\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9461\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44649\
        );

    \I__9460\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44649\
        );

    \I__9459\ : InMux
    port map (
            O => \N__44654\,
            I => \N__44646\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__44649\,
            I => \N__44643\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__44646\,
            I => \N__44640\
        );

    \I__9456\ : Odrv4
    port map (
            O => \N__44643\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__44640\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__9454\ : InMux
    port map (
            O => \N__44635\,
            I => \N__44632\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__44632\,
            I => \N__44629\
        );

    \I__9452\ : Odrv12
    port map (
            O => \N__44629\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__9451\ : CascadeMux
    port map (
            O => \N__44626\,
            I => \N__44623\
        );

    \I__9450\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44620\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__44620\,
            I => \N__44617\
        );

    \I__9448\ : Span4Mux_h
    port map (
            O => \N__44617\,
            I => \N__44614\
        );

    \I__9447\ : Span4Mux_v
    port map (
            O => \N__44614\,
            I => \N__44611\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__44611\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__9445\ : CascadeMux
    port map (
            O => \N__44608\,
            I => \N__44605\
        );

    \I__9444\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44602\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__44602\,
            I => \N__44599\
        );

    \I__9442\ : Span4Mux_h
    port map (
            O => \N__44599\,
            I => \N__44596\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__44596\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__9440\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44590\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__44590\,
            I => \N__44587\
        );

    \I__9438\ : Odrv12
    port map (
            O => \N__44587\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__9437\ : InMux
    port map (
            O => \N__44584\,
            I => \N__44581\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__44581\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__9435\ : InMux
    port map (
            O => \N__44578\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__9434\ : InMux
    port map (
            O => \N__44575\,
            I => \N__44569\
        );

    \I__9433\ : InMux
    port map (
            O => \N__44574\,
            I => \N__44569\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__44569\,
            I => \N__44565\
        );

    \I__9431\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44562\
        );

    \I__9430\ : Span4Mux_v
    port map (
            O => \N__44565\,
            I => \N__44556\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__44562\,
            I => \N__44556\
        );

    \I__9428\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44553\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__44556\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__44553\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__44548\,
            I => \N__44544\
        );

    \I__9424\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44540\
        );

    \I__9423\ : InMux
    port map (
            O => \N__44544\,
            I => \N__44535\
        );

    \I__9422\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44535\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__44540\,
            I => \N__44532\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__44535\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9419\ : Odrv4
    port map (
            O => \N__44532\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9418\ : CascadeMux
    port map (
            O => \N__44527\,
            I => \N__44523\
        );

    \I__9417\ : CascadeMux
    port map (
            O => \N__44526\,
            I => \N__44520\
        );

    \I__9416\ : InMux
    port map (
            O => \N__44523\,
            I => \N__44517\
        );

    \I__9415\ : InMux
    port map (
            O => \N__44520\,
            I => \N__44514\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__44517\,
            I => \N__44510\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__44514\,
            I => \N__44507\
        );

    \I__9412\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44504\
        );

    \I__9411\ : Span4Mux_v
    port map (
            O => \N__44510\,
            I => \N__44498\
        );

    \I__9410\ : Span4Mux_v
    port map (
            O => \N__44507\,
            I => \N__44498\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__44504\,
            I => \N__44495\
        );

    \I__9408\ : InMux
    port map (
            O => \N__44503\,
            I => \N__44492\
        );

    \I__9407\ : Odrv4
    port map (
            O => \N__44498\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9406\ : Odrv4
    port map (
            O => \N__44495\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__44492\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9404\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44481\
        );

    \I__9403\ : InMux
    port map (
            O => \N__44484\,
            I => \N__44478\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44474\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__44478\,
            I => \N__44471\
        );

    \I__9400\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44468\
        );

    \I__9399\ : Odrv12
    port map (
            O => \N__44474\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__44471\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__44468\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9396\ : InMux
    port map (
            O => \N__44461\,
            I => \N__44457\
        );

    \I__9395\ : InMux
    port map (
            O => \N__44460\,
            I => \N__44454\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__44457\,
            I => \N__44450\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__44454\,
            I => \N__44447\
        );

    \I__9392\ : InMux
    port map (
            O => \N__44453\,
            I => \N__44444\
        );

    \I__9391\ : Span4Mux_h
    port map (
            O => \N__44450\,
            I => \N__44440\
        );

    \I__9390\ : Span4Mux_v
    port map (
            O => \N__44447\,
            I => \N__44435\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__44444\,
            I => \N__44435\
        );

    \I__9388\ : InMux
    port map (
            O => \N__44443\,
            I => \N__44432\
        );

    \I__9387\ : Odrv4
    port map (
            O => \N__44440\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9386\ : Odrv4
    port map (
            O => \N__44435\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__44432\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9384\ : CascadeMux
    port map (
            O => \N__44425\,
            I => \N__44422\
        );

    \I__9383\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44418\
        );

    \I__9382\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44415\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__44418\,
            I => \N__44411\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__44415\,
            I => \N__44408\
        );

    \I__9379\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44405\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__44411\,
            I => \N__44398\
        );

    \I__9377\ : Span4Mux_v
    port map (
            O => \N__44408\,
            I => \N__44398\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__44405\,
            I => \N__44398\
        );

    \I__9375\ : Odrv4
    port map (
            O => \N__44398\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9374\ : CascadeMux
    port map (
            O => \N__44395\,
            I => \N__44392\
        );

    \I__9373\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44387\
        );

    \I__9372\ : InMux
    port map (
            O => \N__44391\,
            I => \N__44384\
        );

    \I__9371\ : CascadeMux
    port map (
            O => \N__44390\,
            I => \N__44381\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__44387\,
            I => \N__44378\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__44384\,
            I => \N__44375\
        );

    \I__9368\ : InMux
    port map (
            O => \N__44381\,
            I => \N__44372\
        );

    \I__9367\ : Span4Mux_v
    port map (
            O => \N__44378\,
            I => \N__44366\
        );

    \I__9366\ : Span4Mux_v
    port map (
            O => \N__44375\,
            I => \N__44366\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__44372\,
            I => \N__44363\
        );

    \I__9364\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44360\
        );

    \I__9363\ : Odrv4
    port map (
            O => \N__44366\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9362\ : Odrv12
    port map (
            O => \N__44363\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__44360\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9360\ : InMux
    port map (
            O => \N__44353\,
            I => \N__44350\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__44350\,
            I => \N__44345\
        );

    \I__9358\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44342\
        );

    \I__9357\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44339\
        );

    \I__9356\ : Span4Mux_v
    port map (
            O => \N__44345\,
            I => \N__44334\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__44342\,
            I => \N__44334\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__44339\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9353\ : Odrv4
    port map (
            O => \N__44334\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9352\ : CascadeMux
    port map (
            O => \N__44329\,
            I => \N__44325\
        );

    \I__9351\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44321\
        );

    \I__9350\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44315\
        );

    \I__9349\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44315\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__44321\,
            I => \N__44312\
        );

    \I__9347\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44309\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__44315\,
            I => \N__44306\
        );

    \I__9345\ : Span4Mux_v
    port map (
            O => \N__44312\,
            I => \N__44299\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__44309\,
            I => \N__44299\
        );

    \I__9343\ : Span4Mux_v
    port map (
            O => \N__44306\,
            I => \N__44299\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__44299\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9341\ : InMux
    port map (
            O => \N__44296\,
            I => \N__44293\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44288\
        );

    \I__9339\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44285\
        );

    \I__9338\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44282\
        );

    \I__9337\ : Span4Mux_v
    port map (
            O => \N__44288\,
            I => \N__44277\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__44285\,
            I => \N__44277\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__44282\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__44277\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9333\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44266\
        );

    \I__9332\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44266\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__44266\,
            I => \N__44261\
        );

    \I__9330\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44258\
        );

    \I__9329\ : InMux
    port map (
            O => \N__44264\,
            I => \N__44255\
        );

    \I__9328\ : Odrv12
    port map (
            O => \N__44261\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__44258\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__44255\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9325\ : CascadeMux
    port map (
            O => \N__44248\,
            I => \N__44244\
        );

    \I__9324\ : InMux
    port map (
            O => \N__44247\,
            I => \N__44238\
        );

    \I__9323\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44238\
        );

    \I__9322\ : InMux
    port map (
            O => \N__44243\,
            I => \N__44235\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__44238\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__44235\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9319\ : InMux
    port map (
            O => \N__44230\,
            I => \N__44227\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__44227\,
            I => \N__44223\
        );

    \I__9317\ : InMux
    port map (
            O => \N__44226\,
            I => \N__44220\
        );

    \I__9316\ : Span4Mux_h
    port map (
            O => \N__44223\,
            I => \N__44217\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__44220\,
            I => \N__44214\
        );

    \I__9314\ : Span4Mux_v
    port map (
            O => \N__44217\,
            I => \N__44210\
        );

    \I__9313\ : Span4Mux_v
    port map (
            O => \N__44214\,
            I => \N__44207\
        );

    \I__9312\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44204\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__44210\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9310\ : Odrv4
    port map (
            O => \N__44207\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__44204\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9308\ : CEMux
    port map (
            O => \N__44197\,
            I => \N__44176\
        );

    \I__9307\ : CEMux
    port map (
            O => \N__44196\,
            I => \N__44176\
        );

    \I__9306\ : CEMux
    port map (
            O => \N__44195\,
            I => \N__44176\
        );

    \I__9305\ : CEMux
    port map (
            O => \N__44194\,
            I => \N__44176\
        );

    \I__9304\ : CEMux
    port map (
            O => \N__44193\,
            I => \N__44176\
        );

    \I__9303\ : CEMux
    port map (
            O => \N__44192\,
            I => \N__44176\
        );

    \I__9302\ : CEMux
    port map (
            O => \N__44191\,
            I => \N__44176\
        );

    \I__9301\ : GlobalMux
    port map (
            O => \N__44176\,
            I => \N__44173\
        );

    \I__9300\ : gio2CtrlBuf
    port map (
            O => \N__44173\,
            I => \current_shift_inst.timer_s1.N_163_i_g\
        );

    \I__9299\ : CascadeMux
    port map (
            O => \N__44170\,
            I => \N__44167\
        );

    \I__9298\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44161\
        );

    \I__9297\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44161\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__44161\,
            I => \N__44157\
        );

    \I__9295\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44154\
        );

    \I__9294\ : Odrv4
    port map (
            O => \N__44157\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__44154\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9292\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44144\
        );

    \I__9291\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44139\
        );

    \I__9290\ : InMux
    port map (
            O => \N__44147\,
            I => \N__44139\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__44144\,
            I => \N__44136\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__44139\,
            I => \N__44132\
        );

    \I__9287\ : Span4Mux_v
    port map (
            O => \N__44136\,
            I => \N__44129\
        );

    \I__9286\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44126\
        );

    \I__9285\ : Odrv4
    port map (
            O => \N__44132\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__44129\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__44126\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__9282\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44115\
        );

    \I__9281\ : CascadeMux
    port map (
            O => \N__44118\,
            I => \N__44111\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__44115\,
            I => \N__44108\
        );

    \I__9279\ : InMux
    port map (
            O => \N__44114\,
            I => \N__44105\
        );

    \I__9278\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44102\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__44108\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__44105\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__44102\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__9274\ : InMux
    port map (
            O => \N__44095\,
            I => \N__44092\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__44092\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__44089\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__9271\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44082\
        );

    \I__9270\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44079\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44072\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__44079\,
            I => \N__44072\
        );

    \I__9267\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44067\
        );

    \I__9266\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44067\
        );

    \I__9265\ : Odrv4
    port map (
            O => \N__44072\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__44067\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__9263\ : CascadeMux
    port map (
            O => \N__44062\,
            I => \N__44058\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__44061\,
            I => \N__44055\
        );

    \I__9261\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44052\
        );

    \I__9260\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44049\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44046\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__44039\
        );

    \I__9257\ : Span4Mux_v
    port map (
            O => \N__44046\,
            I => \N__44039\
        );

    \I__9256\ : InMux
    port map (
            O => \N__44045\,
            I => \N__44036\
        );

    \I__9255\ : InMux
    port map (
            O => \N__44044\,
            I => \N__44033\
        );

    \I__9254\ : Odrv4
    port map (
            O => \N__44039\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__44036\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__44033\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9251\ : InMux
    port map (
            O => \N__44026\,
            I => \N__44023\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__44023\,
            I => \N__44018\
        );

    \I__9249\ : InMux
    port map (
            O => \N__44022\,
            I => \N__44015\
        );

    \I__9248\ : InMux
    port map (
            O => \N__44021\,
            I => \N__44012\
        );

    \I__9247\ : Odrv4
    port map (
            O => \N__44018\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__44015\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__44012\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__9244\ : InMux
    port map (
            O => \N__44005\,
            I => \N__44002\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__44002\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9242\ : InMux
    port map (
            O => \N__43999\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9241\ : InMux
    port map (
            O => \N__43996\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9240\ : InMux
    port map (
            O => \N__43993\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9239\ : InMux
    port map (
            O => \N__43990\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9238\ : InMux
    port map (
            O => \N__43987\,
            I => \bfn_17_13_0_\
        );

    \I__9237\ : InMux
    port map (
            O => \N__43984\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9236\ : InMux
    port map (
            O => \N__43981\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9235\ : InMux
    port map (
            O => \N__43978\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9234\ : InMux
    port map (
            O => \N__43975\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9233\ : CEMux
    port map (
            O => \N__43972\,
            I => \N__43967\
        );

    \I__9232\ : CEMux
    port map (
            O => \N__43971\,
            I => \N__43964\
        );

    \I__9231\ : CEMux
    port map (
            O => \N__43970\,
            I => \N__43960\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__43967\,
            I => \N__43956\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__43964\,
            I => \N__43953\
        );

    \I__9228\ : CEMux
    port map (
            O => \N__43963\,
            I => \N__43950\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__43960\,
            I => \N__43947\
        );

    \I__9226\ : CEMux
    port map (
            O => \N__43959\,
            I => \N__43944\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__43956\,
            I => \N__43941\
        );

    \I__9224\ : Span4Mux_h
    port map (
            O => \N__43953\,
            I => \N__43938\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__43950\,
            I => \N__43935\
        );

    \I__9222\ : Span4Mux_h
    port map (
            O => \N__43947\,
            I => \N__43930\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__43944\,
            I => \N__43930\
        );

    \I__9220\ : Span4Mux_h
    port map (
            O => \N__43941\,
            I => \N__43927\
        );

    \I__9219\ : Span4Mux_h
    port map (
            O => \N__43938\,
            I => \N__43924\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__43935\,
            I => \N__43921\
        );

    \I__9217\ : Span4Mux_h
    port map (
            O => \N__43930\,
            I => \N__43918\
        );

    \I__9216\ : Odrv4
    port map (
            O => \N__43927\,
            I => \delay_measurement_inst.delay_hc_timer.N_165_i\
        );

    \I__9215\ : Odrv4
    port map (
            O => \N__43924\,
            I => \delay_measurement_inst.delay_hc_timer.N_165_i\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__43921\,
            I => \delay_measurement_inst.delay_hc_timer.N_165_i\
        );

    \I__9213\ : Odrv4
    port map (
            O => \N__43918\,
            I => \delay_measurement_inst.delay_hc_timer.N_165_i\
        );

    \I__9212\ : InMux
    port map (
            O => \N__43909\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9211\ : InMux
    port map (
            O => \N__43906\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9210\ : InMux
    port map (
            O => \N__43903\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9209\ : InMux
    port map (
            O => \N__43900\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9208\ : InMux
    port map (
            O => \N__43897\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9207\ : InMux
    port map (
            O => \N__43894\,
            I => \bfn_17_12_0_\
        );

    \I__9206\ : InMux
    port map (
            O => \N__43891\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9205\ : InMux
    port map (
            O => \N__43888\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9204\ : InMux
    port map (
            O => \N__43885\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9203\ : InMux
    port map (
            O => \N__43882\,
            I => \N__43879\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__43879\,
            I => \N__43875\
        );

    \I__9201\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43872\
        );

    \I__9200\ : Odrv4
    port map (
            O => \N__43875\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__43872\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__9198\ : InMux
    port map (
            O => \N__43867\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9197\ : InMux
    port map (
            O => \N__43864\,
            I => \N__43860\
        );

    \I__9196\ : InMux
    port map (
            O => \N__43863\,
            I => \N__43857\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__43860\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__43857\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__9193\ : InMux
    port map (
            O => \N__43852\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9192\ : InMux
    port map (
            O => \N__43849\,
            I => \N__43845\
        );

    \I__9191\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43842\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__43845\,
            I => \N__43839\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__43842\,
            I => \N__43836\
        );

    \I__9188\ : Span4Mux_v
    port map (
            O => \N__43839\,
            I => \N__43833\
        );

    \I__9187\ : Odrv12
    port map (
            O => \N__43836\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__43833\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__9185\ : InMux
    port map (
            O => \N__43828\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__43825\,
            I => \N__43822\
        );

    \I__9183\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43818\
        );

    \I__9182\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43815\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__43818\,
            I => \N__43812\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__43815\,
            I => \N__43809\
        );

    \I__9179\ : Span4Mux_v
    port map (
            O => \N__43812\,
            I => \N__43806\
        );

    \I__9178\ : Odrv4
    port map (
            O => \N__43809\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__9177\ : Odrv4
    port map (
            O => \N__43806\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__9176\ : InMux
    port map (
            O => \N__43801\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9175\ : InMux
    port map (
            O => \N__43798\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9174\ : InMux
    port map (
            O => \N__43795\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9173\ : InMux
    port map (
            O => \N__43792\,
            I => \bfn_17_11_0_\
        );

    \I__9172\ : InMux
    port map (
            O => \N__43789\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9171\ : InMux
    port map (
            O => \N__43786\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9170\ : InMux
    port map (
            O => \N__43783\,
            I => \N__43780\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__43780\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__43777\,
            I => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\
        );

    \I__9167\ : InMux
    port map (
            O => \N__43774\,
            I => \N__43771\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__43771\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\
        );

    \I__9165\ : InMux
    port map (
            O => \N__43768\,
            I => \N__43765\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__43765\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__43762\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\
        );

    \I__9162\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43756\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__43756\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\
        );

    \I__9160\ : InMux
    port map (
            O => \N__43753\,
            I => \N__43747\
        );

    \I__9159\ : InMux
    port map (
            O => \N__43752\,
            I => \N__43747\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__43747\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__9157\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43741\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__43741\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\
        );

    \I__9155\ : InMux
    port map (
            O => \N__43738\,
            I => \N__43732\
        );

    \I__9154\ : InMux
    port map (
            O => \N__43737\,
            I => \N__43732\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__43732\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__9152\ : InMux
    port map (
            O => \N__43729\,
            I => \N__43726\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__43726\,
            I => \N__43722\
        );

    \I__9150\ : InMux
    port map (
            O => \N__43725\,
            I => \N__43719\
        );

    \I__9149\ : Span4Mux_v
    port map (
            O => \N__43722\,
            I => \N__43714\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__43719\,
            I => \N__43714\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__43714\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9146\ : InMux
    port map (
            O => \N__43711\,
            I => \N__43707\
        );

    \I__9145\ : CascadeMux
    port map (
            O => \N__43710\,
            I => \N__43704\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__43707\,
            I => \N__43701\
        );

    \I__9143\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43698\
        );

    \I__9142\ : Span4Mux_v
    port map (
            O => \N__43701\,
            I => \N__43693\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__43698\,
            I => \N__43693\
        );

    \I__9140\ : Odrv4
    port map (
            O => \N__43693\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__9139\ : InMux
    port map (
            O => \N__43690\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9138\ : InMux
    port map (
            O => \N__43687\,
            I => \N__43684\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__43684\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__9136\ : CascadeMux
    port map (
            O => \N__43681\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\
        );

    \I__9135\ : InMux
    port map (
            O => \N__43678\,
            I => \N__43675\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__43675\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\
        );

    \I__9133\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43669\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__43669\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__43666\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\
        );

    \I__9130\ : InMux
    port map (
            O => \N__43663\,
            I => \N__43660\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__43660\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\
        );

    \I__9128\ : InMux
    port map (
            O => \N__43657\,
            I => \N__43651\
        );

    \I__9127\ : InMux
    port map (
            O => \N__43656\,
            I => \N__43651\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__43651\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__9125\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43645\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__43645\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\
        );

    \I__9123\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43639\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__43639\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__43636\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\
        );

    \I__9120\ : InMux
    port map (
            O => \N__43633\,
            I => \N__43630\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__43630\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\
        );

    \I__9118\ : InMux
    port map (
            O => \N__43627\,
            I => \N__43624\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__43624\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\
        );

    \I__9116\ : InMux
    port map (
            O => \N__43621\,
            I => \N__43616\
        );

    \I__9115\ : InMux
    port map (
            O => \N__43620\,
            I => \N__43613\
        );

    \I__9114\ : InMux
    port map (
            O => \N__43619\,
            I => \N__43610\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__43616\,
            I => \N__43605\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43605\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__43610\,
            I => \N__43602\
        );

    \I__9110\ : Odrv12
    port map (
            O => \N__43605\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9109\ : Odrv4
    port map (
            O => \N__43602\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9108\ : InMux
    port map (
            O => \N__43597\,
            I => \N__43594\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__43594\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__9106\ : CascadeMux
    port map (
            O => \N__43591\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\
        );

    \I__9105\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43585\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__43585\,
            I => \N__43582\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__43582\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\
        );

    \I__9102\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43575\
        );

    \I__9101\ : InMux
    port map (
            O => \N__43578\,
            I => \N__43572\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__43575\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__43572\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__9098\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43564\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__43564\,
            I => \N__43561\
        );

    \I__9096\ : Span4Mux_v
    port map (
            O => \N__43561\,
            I => \N__43558\
        );

    \I__9095\ : Odrv4
    port map (
            O => \N__43558\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\
        );

    \I__9094\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43552\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__43552\,
            I => \N__43549\
        );

    \I__9092\ : Span4Mux_v
    port map (
            O => \N__43549\,
            I => \N__43546\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__43546\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\
        );

    \I__9090\ : InMux
    port map (
            O => \N__43543\,
            I => \N__43540\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__43540\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__9088\ : CascadeMux
    port map (
            O => \N__43537\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\
        );

    \I__9087\ : InMux
    port map (
            O => \N__43534\,
            I => \N__43531\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__43531\,
            I => \N__43528\
        );

    \I__9085\ : Odrv4
    port map (
            O => \N__43528\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\
        );

    \I__9084\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43522\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__43522\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__9082\ : CascadeMux
    port map (
            O => \N__43519\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\
        );

    \I__9081\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43513\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__43513\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\
        );

    \I__9079\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43507\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__43507\,
            I => \N__43504\
        );

    \I__9077\ : Odrv4
    port map (
            O => \N__43504\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__9076\ : CascadeMux
    port map (
            O => \N__43501\,
            I => \N__43497\
        );

    \I__9075\ : InMux
    port map (
            O => \N__43500\,
            I => \N__43494\
        );

    \I__9074\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43491\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__43494\,
            I => \N__43484\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__43491\,
            I => \N__43484\
        );

    \I__9071\ : InMux
    port map (
            O => \N__43490\,
            I => \N__43481\
        );

    \I__9070\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43478\
        );

    \I__9069\ : Span4Mux_v
    port map (
            O => \N__43484\,
            I => \N__43471\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__43481\,
            I => \N__43471\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__43478\,
            I => \N__43471\
        );

    \I__9066\ : Odrv4
    port map (
            O => \N__43471\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9065\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43464\
        );

    \I__9064\ : InMux
    port map (
            O => \N__43467\,
            I => \N__43461\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__43464\,
            I => \N__43457\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__43461\,
            I => \N__43454\
        );

    \I__9061\ : InMux
    port map (
            O => \N__43460\,
            I => \N__43451\
        );

    \I__9060\ : Span4Mux_v
    port map (
            O => \N__43457\,
            I => \N__43448\
        );

    \I__9059\ : Span4Mux_v
    port map (
            O => \N__43454\,
            I => \N__43443\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__43451\,
            I => \N__43443\
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__43448\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9056\ : Odrv4
    port map (
            O => \N__43443\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9055\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43435\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__43435\,
            I => \N__43432\
        );

    \I__9053\ : Odrv12
    port map (
            O => \N__43432\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__9052\ : InMux
    port map (
            O => \N__43429\,
            I => \N__43426\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__43426\,
            I => \N__43423\
        );

    \I__9050\ : Odrv4
    port map (
            O => \N__43423\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__9049\ : CascadeMux
    port map (
            O => \N__43420\,
            I => \N__43416\
        );

    \I__9048\ : CascadeMux
    port map (
            O => \N__43419\,
            I => \N__43413\
        );

    \I__9047\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43410\
        );

    \I__9046\ : InMux
    port map (
            O => \N__43413\,
            I => \N__43407\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__43410\,
            I => \N__43403\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__43407\,
            I => \N__43400\
        );

    \I__9043\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43397\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__43403\,
            I => \N__43389\
        );

    \I__9041\ : Span4Mux_v
    port map (
            O => \N__43400\,
            I => \N__43389\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__43397\,
            I => \N__43389\
        );

    \I__9039\ : InMux
    port map (
            O => \N__43396\,
            I => \N__43386\
        );

    \I__9038\ : Odrv4
    port map (
            O => \N__43389\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__43386\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9036\ : InMux
    port map (
            O => \N__43381\,
            I => \N__43376\
        );

    \I__9035\ : InMux
    port map (
            O => \N__43380\,
            I => \N__43373\
        );

    \I__9034\ : InMux
    port map (
            O => \N__43379\,
            I => \N__43370\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__43376\,
            I => \N__43365\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__43373\,
            I => \N__43365\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__43370\,
            I => \N__43362\
        );

    \I__9030\ : Odrv12
    port map (
            O => \N__43365\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__43362\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9028\ : InMux
    port map (
            O => \N__43357\,
            I => \N__43354\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__43354\,
            I => \N__43351\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__43351\,
            I => \N__43348\
        );

    \I__9025\ : Odrv4
    port map (
            O => \N__43348\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__9024\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43342\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__43342\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__9022\ : CascadeMux
    port map (
            O => \N__43339\,
            I => \N__43336\
        );

    \I__9021\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43333\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43330\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__43330\,
            I => \N__43327\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__43327\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__9017\ : InMux
    port map (
            O => \N__43324\,
            I => \N__43321\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__43321\,
            I => \N__43318\
        );

    \I__9015\ : Span4Mux_h
    port map (
            O => \N__43318\,
            I => \N__43315\
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__43315\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__9013\ : InMux
    port map (
            O => \N__43312\,
            I => \N__43309\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__43309\,
            I => \N__43306\
        );

    \I__9011\ : Span4Mux_h
    port map (
            O => \N__43306\,
            I => \N__43303\
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__43303\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__9009\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43297\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43294\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__43294\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__9006\ : InMux
    port map (
            O => \N__43291\,
            I => \N__43288\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__43288\,
            I => \N__43285\
        );

    \I__9004\ : Odrv4
    port map (
            O => \N__43285\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__9003\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43279\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__43279\,
            I => \N__43276\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__43276\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__9000\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43270\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__43270\,
            I => \N__43267\
        );

    \I__8998\ : Odrv4
    port map (
            O => \N__43267\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__8997\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43261\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__43261\,
            I => \N__43258\
        );

    \I__8995\ : Span4Mux_h
    port map (
            O => \N__43258\,
            I => \N__43255\
        );

    \I__8994\ : Odrv4
    port map (
            O => \N__43255\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__8993\ : InMux
    port map (
            O => \N__43252\,
            I => \N__43249\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__43249\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8991\ : InMux
    port map (
            O => \N__43246\,
            I => \N__43243\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__43243\,
            I => \N__43240\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__43240\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__8988\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43224\
        );

    \I__8987\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43224\
        );

    \I__8986\ : InMux
    port map (
            O => \N__43235\,
            I => \N__43207\
        );

    \I__8985\ : InMux
    port map (
            O => \N__43234\,
            I => \N__43207\
        );

    \I__8984\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43207\
        );

    \I__8983\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43207\
        );

    \I__8982\ : InMux
    port map (
            O => \N__43231\,
            I => \N__43207\
        );

    \I__8981\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43202\
        );

    \I__8980\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43202\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__43224\,
            I => \N__43199\
        );

    \I__8978\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43192\
        );

    \I__8977\ : InMux
    port map (
            O => \N__43222\,
            I => \N__43192\
        );

    \I__8976\ : InMux
    port map (
            O => \N__43221\,
            I => \N__43192\
        );

    \I__8975\ : InMux
    port map (
            O => \N__43220\,
            I => \N__43185\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43185\
        );

    \I__8973\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43185\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__43207\,
            I => \N__43170\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__43202\,
            I => \N__43170\
        );

    \I__8970\ : Span4Mux_v
    port map (
            O => \N__43199\,
            I => \N__43163\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__43192\,
            I => \N__43163\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__43185\,
            I => \N__43163\
        );

    \I__8967\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43154\
        );

    \I__8966\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43154\
        );

    \I__8965\ : InMux
    port map (
            O => \N__43182\,
            I => \N__43154\
        );

    \I__8964\ : InMux
    port map (
            O => \N__43181\,
            I => \N__43154\
        );

    \I__8963\ : InMux
    port map (
            O => \N__43180\,
            I => \N__43147\
        );

    \I__8962\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43147\
        );

    \I__8961\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43147\
        );

    \I__8960\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43144\
        );

    \I__8959\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43139\
        );

    \I__8958\ : InMux
    port map (
            O => \N__43175\,
            I => \N__43139\
        );

    \I__8957\ : Odrv12
    port map (
            O => \N__43170\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8956\ : Odrv4
    port map (
            O => \N__43163\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__43154\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__43147\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__43144\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__43139\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__43126\,
            I => \N__43123\
        );

    \I__8950\ : InMux
    port map (
            O => \N__43123\,
            I => \N__43120\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__43120\,
            I => \N__43117\
        );

    \I__8948\ : Odrv4
    port map (
            O => \N__43117\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__8947\ : InMux
    port map (
            O => \N__43114\,
            I => \N__43111\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__43111\,
            I => \N__43108\
        );

    \I__8945\ : Span4Mux_h
    port map (
            O => \N__43108\,
            I => \N__43105\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__43105\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__8943\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43099\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__43099\,
            I => \N__43096\
        );

    \I__8941\ : Odrv4
    port map (
            O => \N__43096\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__8940\ : CascadeMux
    port map (
            O => \N__43093\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__8939\ : CascadeMux
    port map (
            O => \N__43090\,
            I => \N__43086\
        );

    \I__8938\ : InMux
    port map (
            O => \N__43089\,
            I => \N__43082\
        );

    \I__8937\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43079\
        );

    \I__8936\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43076\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43071\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__43079\,
            I => \N__43071\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__43076\,
            I => \current_shift_inst.N_1379_i\
        );

    \I__8932\ : Odrv4
    port map (
            O => \N__43071\,
            I => \current_shift_inst.N_1379_i\
        );

    \I__8931\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43063\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__43063\,
            I => \N__43060\
        );

    \I__8929\ : Span4Mux_h
    port map (
            O => \N__43060\,
            I => \N__43057\
        );

    \I__8928\ : Odrv4
    port map (
            O => \N__43057\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__43054\,
            I => \N__43051\
        );

    \I__8926\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43048\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__43048\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8924\ : InMux
    port map (
            O => \N__43045\,
            I => \N__43042\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__43042\,
            I => \N__43039\
        );

    \I__8922\ : Odrv4
    port map (
            O => \N__43039\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__8921\ : CascadeMux
    port map (
            O => \N__43036\,
            I => \N__43033\
        );

    \I__8920\ : InMux
    port map (
            O => \N__43033\,
            I => \N__43030\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__43030\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8918\ : CascadeMux
    port map (
            O => \N__43027\,
            I => \N__43024\
        );

    \I__8917\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43021\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__43021\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__43018\,
            I => \N__43015\
        );

    \I__8914\ : InMux
    port map (
            O => \N__43015\,
            I => \N__43012\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__43012\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__8912\ : InMux
    port map (
            O => \N__43009\,
            I => \N__43006\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__43006\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__8910\ : CascadeMux
    port map (
            O => \N__43003\,
            I => \N__43000\
        );

    \I__8909\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42997\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__42997\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8907\ : CascadeMux
    port map (
            O => \N__42994\,
            I => \N__42991\
        );

    \I__8906\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42988\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__42988\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__8904\ : CascadeMux
    port map (
            O => \N__42985\,
            I => \N__42982\
        );

    \I__8903\ : InMux
    port map (
            O => \N__42982\,
            I => \N__42979\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__42979\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__8901\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42973\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__42973\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__8899\ : InMux
    port map (
            O => \N__42970\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__8898\ : InMux
    port map (
            O => \N__42967\,
            I => \N__42964\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__42964\,
            I => \N__42961\
        );

    \I__8896\ : Span4Mux_h
    port map (
            O => \N__42961\,
            I => \N__42958\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__42958\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__8894\ : InMux
    port map (
            O => \N__42955\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__8893\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42949\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__42949\,
            I => \N__42946\
        );

    \I__8891\ : Span4Mux_h
    port map (
            O => \N__42946\,
            I => \N__42943\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__42943\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__8889\ : InMux
    port map (
            O => \N__42940\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__8888\ : InMux
    port map (
            O => \N__42937\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__8887\ : InMux
    port map (
            O => \N__42934\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__8886\ : InMux
    port map (
            O => \N__42931\,
            I => \N__42928\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__42928\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__8884\ : CascadeMux
    port map (
            O => \N__42925\,
            I => \N__42922\
        );

    \I__8883\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42919\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__42919\,
            I => \N__42916\
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__42916\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__8880\ : CascadeMux
    port map (
            O => \N__42913\,
            I => \N__42910\
        );

    \I__8879\ : InMux
    port map (
            O => \N__42910\,
            I => \N__42907\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__42907\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__8877\ : InMux
    port map (
            O => \N__42904\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__8876\ : InMux
    port map (
            O => \N__42901\,
            I => \N__42898\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__8874\ : Odrv12
    port map (
            O => \N__42895\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__8873\ : InMux
    port map (
            O => \N__42892\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__8872\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42886\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__42886\,
            I => \N__42883\
        );

    \I__8870\ : Span4Mux_h
    port map (
            O => \N__42883\,
            I => \N__42880\
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__42880\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__8868\ : InMux
    port map (
            O => \N__42877\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__8867\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42871\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42868\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__42868\,
            I => \N__42865\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__42865\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__8863\ : InMux
    port map (
            O => \N__42862\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__8862\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42856\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__42856\,
            I => \N__42853\
        );

    \I__8860\ : Span4Mux_h
    port map (
            O => \N__42853\,
            I => \N__42850\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__42850\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__8858\ : InMux
    port map (
            O => \N__42847\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__8857\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42841\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__42841\,
            I => \N__42838\
        );

    \I__8855\ : Span4Mux_h
    port map (
            O => \N__42838\,
            I => \N__42835\
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__42835\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__8853\ : InMux
    port map (
            O => \N__42832\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__8852\ : InMux
    port map (
            O => \N__42829\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__8851\ : InMux
    port map (
            O => \N__42826\,
            I => \bfn_16_16_0_\
        );

    \I__8850\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42820\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__42820\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__8848\ : InMux
    port map (
            O => \N__42817\,
            I => \bfn_16_14_0_\
        );

    \I__8847\ : InMux
    port map (
            O => \N__42814\,
            I => \N__42811\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__42811\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__8845\ : InMux
    port map (
            O => \N__42808\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__8844\ : InMux
    port map (
            O => \N__42805\,
            I => \N__42802\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__42802\,
            I => \N__42799\
        );

    \I__8842\ : Span4Mux_h
    port map (
            O => \N__42799\,
            I => \N__42796\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__42796\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__8840\ : InMux
    port map (
            O => \N__42793\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__8839\ : InMux
    port map (
            O => \N__42790\,
            I => \N__42787\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__42787\,
            I => \N__42784\
        );

    \I__8837\ : Span4Mux_v
    port map (
            O => \N__42784\,
            I => \N__42781\
        );

    \I__8836\ : Odrv4
    port map (
            O => \N__42781\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__8835\ : InMux
    port map (
            O => \N__42778\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__8834\ : InMux
    port map (
            O => \N__42775\,
            I => \N__42772\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__42772\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__8832\ : InMux
    port map (
            O => \N__42769\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__8831\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42763\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__42763\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__8829\ : InMux
    port map (
            O => \N__42760\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__8828\ : InMux
    port map (
            O => \N__42757\,
            I => \N__42754\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__42754\,
            I => \N__42751\
        );

    \I__8826\ : Span4Mux_h
    port map (
            O => \N__42751\,
            I => \N__42748\
        );

    \I__8825\ : Odrv4
    port map (
            O => \N__42748\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__8824\ : InMux
    port map (
            O => \N__42745\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__8823\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42739\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__42739\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__8821\ : InMux
    port map (
            O => \N__42736\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__8820\ : InMux
    port map (
            O => \N__42733\,
            I => \N__42730\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__42730\,
            I => \N__42727\
        );

    \I__8818\ : Odrv12
    port map (
            O => \N__42727\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__8817\ : InMux
    port map (
            O => \N__42724\,
            I => \bfn_16_15_0_\
        );

    \I__8816\ : InMux
    port map (
            O => \N__42721\,
            I => \N__42718\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__42718\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__8814\ : InMux
    port map (
            O => \N__42715\,
            I => \N__42712\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__42712\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__8812\ : InMux
    port map (
            O => \N__42709\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__8811\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42703\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__42703\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__8809\ : InMux
    port map (
            O => \N__42700\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__8808\ : InMux
    port map (
            O => \N__42697\,
            I => \N__42694\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__42694\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__8806\ : InMux
    port map (
            O => \N__42691\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__8805\ : InMux
    port map (
            O => \N__42688\,
            I => \N__42685\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__42685\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__8803\ : InMux
    port map (
            O => \N__42682\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__8802\ : InMux
    port map (
            O => \N__42679\,
            I => \N__42676\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__42676\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__8800\ : InMux
    port map (
            O => \N__42673\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__8799\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42667\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__42667\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__8797\ : InMux
    port map (
            O => \N__42664\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__8796\ : InMux
    port map (
            O => \N__42661\,
            I => \N__42658\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42655\
        );

    \I__8794\ : Span4Mux_h
    port map (
            O => \N__42655\,
            I => \N__42652\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__42652\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__8792\ : InMux
    port map (
            O => \N__42649\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__8791\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42643\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__42643\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\
        );

    \I__8789\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42636\
        );

    \I__8788\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42632\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__42636\,
            I => \N__42627\
        );

    \I__8786\ : InMux
    port map (
            O => \N__42635\,
            I => \N__42624\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__42632\,
            I => \N__42621\
        );

    \I__8784\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42618\
        );

    \I__8783\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42615\
        );

    \I__8782\ : Odrv4
    port map (
            O => \N__42627\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__42624\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8780\ : Odrv12
    port map (
            O => \N__42621\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__42618\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__42615\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__8777\ : InMux
    port map (
            O => \N__42604\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\
        );

    \I__8776\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42598\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42594\
        );

    \I__8774\ : InMux
    port map (
            O => \N__42597\,
            I => \N__42591\
        );

    \I__8773\ : Span4Mux_h
    port map (
            O => \N__42594\,
            I => \N__42588\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__42591\,
            I => \N__42585\
        );

    \I__8771\ : Odrv4
    port map (
            O => \N__42588\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_28
        );

    \I__8770\ : Odrv12
    port map (
            O => \N__42585\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_28
        );

    \I__8769\ : InMux
    port map (
            O => \N__42580\,
            I => \N__42577\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__42577\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__42574\,
            I => \N__42571\
        );

    \I__8766\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42568\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__42568\,
            I => \N__42565\
        );

    \I__8764\ : Span4Mux_v
    port map (
            O => \N__42565\,
            I => \N__42562\
        );

    \I__8763\ : Odrv4
    port map (
            O => \N__42562\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__42559\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__8761\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42552\
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__42555\,
            I => \N__42549\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42546\
        );

    \I__8758\ : InMux
    port map (
            O => \N__42549\,
            I => \N__42543\
        );

    \I__8757\ : Span4Mux_v
    port map (
            O => \N__42546\,
            I => \N__42540\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__42543\,
            I => \N__42537\
        );

    \I__8755\ : Span4Mux_h
    port map (
            O => \N__42540\,
            I => \N__42532\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__42537\,
            I => \N__42532\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__42532\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__8752\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42526\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__42526\,
            I => \N__42522\
        );

    \I__8750\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42518\
        );

    \I__8749\ : Span4Mux_h
    port map (
            O => \N__42522\,
            I => \N__42515\
        );

    \I__8748\ : InMux
    port map (
            O => \N__42521\,
            I => \N__42512\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__42518\,
            I => \N__42509\
        );

    \I__8746\ : Odrv4
    port map (
            O => \N__42515\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__42512\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8744\ : Odrv12
    port map (
            O => \N__42509\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__8743\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42499\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__42499\,
            I => \N__42495\
        );

    \I__8741\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42492\
        );

    \I__8740\ : Odrv4
    port map (
            O => \N__42495\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__42492\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\
        );

    \I__8738\ : InMux
    port map (
            O => \N__42487\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\
        );

    \I__8737\ : InMux
    port map (
            O => \N__42484\,
            I => \N__42480\
        );

    \I__8736\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42477\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__42480\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__42477\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\
        );

    \I__8733\ : InMux
    port map (
            O => \N__42472\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\
        );

    \I__8732\ : InMux
    port map (
            O => \N__42469\,
            I => \N__42466\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__42466\,
            I => \N__42463\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__42463\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\
        );

    \I__8729\ : InMux
    port map (
            O => \N__42460\,
            I => \N__42456\
        );

    \I__8728\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42453\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__42456\,
            I => \N__42450\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__42453\,
            I => \N__42447\
        );

    \I__8725\ : Odrv4
    port map (
            O => \N__42450\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__42447\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\
        );

    \I__8723\ : InMux
    port map (
            O => \N__42442\,
            I => \bfn_16_11_0_\
        );

    \I__8722\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42435\
        );

    \I__8721\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42432\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__42435\,
            I => \N__42427\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__42432\,
            I => \N__42427\
        );

    \I__8718\ : Odrv4
    port map (
            O => \N__42427\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\
        );

    \I__8717\ : InMux
    port map (
            O => \N__42424\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\
        );

    \I__8716\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42417\
        );

    \I__8715\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42414\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__42417\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__42414\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\
        );

    \I__8712\ : InMux
    port map (
            O => \N__42409\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\
        );

    \I__8711\ : InMux
    port map (
            O => \N__42406\,
            I => \N__42402\
        );

    \I__8710\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42399\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__42402\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__42399\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\
        );

    \I__8707\ : InMux
    port map (
            O => \N__42394\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\
        );

    \I__8706\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42388\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__42388\,
            I => \N__42385\
        );

    \I__8704\ : Odrv12
    port map (
            O => \N__42385\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\
        );

    \I__8703\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42378\
        );

    \I__8702\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42375\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__42378\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__42375\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\
        );

    \I__8699\ : InMux
    port map (
            O => \N__42370\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\
        );

    \I__8698\ : InMux
    port map (
            O => \N__42367\,
            I => \N__42364\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__42364\,
            I => \N__42361\
        );

    \I__8696\ : Span4Mux_h
    port map (
            O => \N__42361\,
            I => \N__42358\
        );

    \I__8695\ : Odrv4
    port map (
            O => \N__42358\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\
        );

    \I__8694\ : InMux
    port map (
            O => \N__42355\,
            I => \N__42351\
        );

    \I__8693\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42348\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__42351\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__42348\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\
        );

    \I__8690\ : InMux
    port map (
            O => \N__42343\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\
        );

    \I__8689\ : InMux
    port map (
            O => \N__42340\,
            I => \N__42336\
        );

    \I__8688\ : InMux
    port map (
            O => \N__42339\,
            I => \N__42333\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__42336\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__42333\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\
        );

    \I__8685\ : InMux
    port map (
            O => \N__42328\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\
        );

    \I__8684\ : InMux
    port map (
            O => \N__42325\,
            I => \N__42321\
        );

    \I__8683\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42318\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__42321\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__42318\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\
        );

    \I__8680\ : InMux
    port map (
            O => \N__42313\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\
        );

    \I__8679\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42306\
        );

    \I__8678\ : InMux
    port map (
            O => \N__42309\,
            I => \N__42303\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__42306\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__42303\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\
        );

    \I__8675\ : InMux
    port map (
            O => \N__42298\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\
        );

    \I__8674\ : InMux
    port map (
            O => \N__42295\,
            I => \N__42291\
        );

    \I__8673\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42288\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__42291\,
            I => \N__42285\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__42288\,
            I => \N__42282\
        );

    \I__8670\ : Odrv4
    port map (
            O => \N__42285\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\
        );

    \I__8669\ : Odrv4
    port map (
            O => \N__42282\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\
        );

    \I__8668\ : InMux
    port map (
            O => \N__42277\,
            I => \bfn_16_10_0_\
        );

    \I__8667\ : InMux
    port map (
            O => \N__42274\,
            I => \N__42270\
        );

    \I__8666\ : InMux
    port map (
            O => \N__42273\,
            I => \N__42267\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__42270\,
            I => \N__42262\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__42267\,
            I => \N__42262\
        );

    \I__8663\ : Odrv4
    port map (
            O => \N__42262\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\
        );

    \I__8662\ : InMux
    port map (
            O => \N__42259\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\
        );

    \I__8661\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42252\
        );

    \I__8660\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42249\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__42252\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__42249\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\
        );

    \I__8657\ : InMux
    port map (
            O => \N__42244\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\
        );

    \I__8656\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42237\
        );

    \I__8655\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42234\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__42237\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__42234\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\
        );

    \I__8652\ : InMux
    port map (
            O => \N__42229\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\
        );

    \I__8651\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42223\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__42223\,
            I => \N__42220\
        );

    \I__8649\ : Span4Mux_h
    port map (
            O => \N__42220\,
            I => \N__42216\
        );

    \I__8648\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42213\
        );

    \I__8647\ : Span4Mux_h
    port map (
            O => \N__42216\,
            I => \N__42210\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__42213\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\
        );

    \I__8645\ : Odrv4
    port map (
            O => \N__42210\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\
        );

    \I__8644\ : InMux
    port map (
            O => \N__42205\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\
        );

    \I__8643\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42199\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__42199\,
            I => \N__42196\
        );

    \I__8641\ : Span4Mux_h
    port map (
            O => \N__42196\,
            I => \N__42193\
        );

    \I__8640\ : Odrv4
    port map (
            O => \N__42193\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\
        );

    \I__8639\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42186\
        );

    \I__8638\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42183\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__42186\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__42183\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\
        );

    \I__8635\ : InMux
    port map (
            O => \N__42178\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\
        );

    \I__8634\ : InMux
    port map (
            O => \N__42175\,
            I => \N__42171\
        );

    \I__8633\ : InMux
    port map (
            O => \N__42174\,
            I => \N__42168\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__42171\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__42168\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\
        );

    \I__8630\ : InMux
    port map (
            O => \N__42163\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\
        );

    \I__8629\ : InMux
    port map (
            O => \N__42160\,
            I => \N__42156\
        );

    \I__8628\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42153\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__42156\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__42153\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\
        );

    \I__8625\ : InMux
    port map (
            O => \N__42148\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\
        );

    \I__8624\ : InMux
    port map (
            O => \N__42145\,
            I => \N__42141\
        );

    \I__8623\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42138\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__42141\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__42138\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\
        );

    \I__8620\ : InMux
    port map (
            O => \N__42133\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\
        );

    \I__8619\ : InMux
    port map (
            O => \N__42130\,
            I => \N__42126\
        );

    \I__8618\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42123\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__42126\,
            I => \N__42120\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__42123\,
            I => \N__42117\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__42120\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__42117\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\
        );

    \I__8613\ : InMux
    port map (
            O => \N__42112\,
            I => \bfn_16_9_0_\
        );

    \I__8612\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42105\
        );

    \I__8611\ : InMux
    port map (
            O => \N__42108\,
            I => \N__42102\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__42105\,
            I => \N__42097\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__42097\
        );

    \I__8608\ : Span4Mux_v
    port map (
            O => \N__42097\,
            I => \N__42094\
        );

    \I__8607\ : Odrv4
    port map (
            O => \N__42094\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\
        );

    \I__8606\ : InMux
    port map (
            O => \N__42091\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\
        );

    \I__8605\ : InMux
    port map (
            O => \N__42088\,
            I => \N__42084\
        );

    \I__8604\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42081\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__42084\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__42081\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\
        );

    \I__8601\ : InMux
    port map (
            O => \N__42076\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\
        );

    \I__8600\ : InMux
    port map (
            O => \N__42073\,
            I => \N__42069\
        );

    \I__8599\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42066\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__42069\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__42066\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\
        );

    \I__8596\ : InMux
    port map (
            O => \N__42061\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\
        );

    \I__8595\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42054\
        );

    \I__8594\ : InMux
    port map (
            O => \N__42057\,
            I => \N__42051\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__42054\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__42051\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\
        );

    \I__8591\ : InMux
    port map (
            O => \N__42046\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\
        );

    \I__8590\ : CEMux
    port map (
            O => \N__42043\,
            I => \N__42040\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__42040\,
            I => \N__42034\
        );

    \I__8588\ : CEMux
    port map (
            O => \N__42039\,
            I => \N__42029\
        );

    \I__8587\ : CEMux
    port map (
            O => \N__42038\,
            I => \N__42026\
        );

    \I__8586\ : CEMux
    port map (
            O => \N__42037\,
            I => \N__42023\
        );

    \I__8585\ : Span4Mux_h
    port map (
            O => \N__42034\,
            I => \N__42019\
        );

    \I__8584\ : CEMux
    port map (
            O => \N__42033\,
            I => \N__42016\
        );

    \I__8583\ : CEMux
    port map (
            O => \N__42032\,
            I => \N__42013\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__42029\,
            I => \N__42010\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__42026\,
            I => \N__42007\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42004\
        );

    \I__8579\ : CEMux
    port map (
            O => \N__42022\,
            I => \N__42001\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__42019\,
            I => \N__41996\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__42016\,
            I => \N__41996\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__42013\,
            I => \N__41993\
        );

    \I__8575\ : Span4Mux_h
    port map (
            O => \N__42010\,
            I => \N__41990\
        );

    \I__8574\ : Span4Mux_h
    port map (
            O => \N__42007\,
            I => \N__41983\
        );

    \I__8573\ : Span4Mux_v
    port map (
            O => \N__42004\,
            I => \N__41983\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__42001\,
            I => \N__41983\
        );

    \I__8571\ : Span4Mux_h
    port map (
            O => \N__41996\,
            I => \N__41978\
        );

    \I__8570\ : Span4Mux_h
    port map (
            O => \N__41993\,
            I => \N__41978\
        );

    \I__8569\ : Span4Mux_v
    port map (
            O => \N__41990\,
            I => \N__41973\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__41983\,
            I => \N__41973\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__41978\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__41973\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__41968\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31_cascade_\
        );

    \I__8564\ : InMux
    port map (
            O => \N__41965\,
            I => \N__41962\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__41962\,
            I => \N__41959\
        );

    \I__8562\ : Span12Mux_s6_v
    port map (
            O => \N__41959\,
            I => \N__41956\
        );

    \I__8561\ : Odrv12
    port map (
            O => \N__41956\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\
        );

    \I__8560\ : CEMux
    port map (
            O => \N__41953\,
            I => \N__41949\
        );

    \I__8559\ : CEMux
    port map (
            O => \N__41952\,
            I => \N__41944\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__41949\,
            I => \N__41941\
        );

    \I__8557\ : CEMux
    port map (
            O => \N__41948\,
            I => \N__41938\
        );

    \I__8556\ : CEMux
    port map (
            O => \N__41947\,
            I => \N__41935\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__41944\,
            I => \N__41929\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__41941\,
            I => \N__41922\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__41938\,
            I => \N__41922\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__41935\,
            I => \N__41922\
        );

    \I__8551\ : CEMux
    port map (
            O => \N__41934\,
            I => \N__41919\
        );

    \I__8550\ : CEMux
    port map (
            O => \N__41933\,
            I => \N__41916\
        );

    \I__8549\ : CEMux
    port map (
            O => \N__41932\,
            I => \N__41912\
        );

    \I__8548\ : Span4Mux_h
    port map (
            O => \N__41929\,
            I => \N__41905\
        );

    \I__8547\ : Span4Mux_v
    port map (
            O => \N__41922\,
            I => \N__41905\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__41919\,
            I => \N__41905\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41902\
        );

    \I__8544\ : CEMux
    port map (
            O => \N__41915\,
            I => \N__41899\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__41912\,
            I => \N__41896\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__41905\,
            I => \N__41893\
        );

    \I__8541\ : Span4Mux_h
    port map (
            O => \N__41902\,
            I => \N__41890\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__41899\,
            I => \N__41887\
        );

    \I__8539\ : Span4Mux_h
    port map (
            O => \N__41896\,
            I => \N__41884\
        );

    \I__8538\ : Odrv4
    port map (
            O => \N__41893\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__8537\ : Odrv4
    port map (
            O => \N__41890\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__8536\ : Odrv4
    port map (
            O => \N__41887\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__41884\,
            I => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\
        );

    \I__8534\ : CascadeMux
    port map (
            O => \N__41875\,
            I => \N__41872\
        );

    \I__8533\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41869\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__41869\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\
        );

    \I__8531\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41863\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__41863\,
            I => \N__41859\
        );

    \I__8529\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41856\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__41859\,
            I => \N__41853\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__41856\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__41853\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__8525\ : InMux
    port map (
            O => \N__41848\,
            I => \N__41845\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__41845\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\
        );

    \I__8523\ : InMux
    port map (
            O => \N__41842\,
            I => \N__41839\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__41839\,
            I => \N__41836\
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__41836\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\
        );

    \I__8520\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41828\
        );

    \I__8519\ : CascadeMux
    port map (
            O => \N__41832\,
            I => \N__41825\
        );

    \I__8518\ : InMux
    port map (
            O => \N__41831\,
            I => \N__41822\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__41828\,
            I => \N__41819\
        );

    \I__8516\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41816\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__41822\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__41819\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__41816\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\
        );

    \I__8512\ : InMux
    port map (
            O => \N__41809\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\
        );

    \I__8511\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41803\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__41803\,
            I => \N__41800\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__41800\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\
        );

    \I__8508\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41793\
        );

    \I__8507\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41790\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__41793\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__41790\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\
        );

    \I__8504\ : InMux
    port map (
            O => \N__41785\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\
        );

    \I__8503\ : InMux
    port map (
            O => \N__41782\,
            I => \N__41778\
        );

    \I__8502\ : InMux
    port map (
            O => \N__41781\,
            I => \N__41775\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__41778\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__41775\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\
        );

    \I__8499\ : InMux
    port map (
            O => \N__41770\,
            I => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\
        );

    \I__8498\ : InMux
    port map (
            O => \N__41767\,
            I => \N__41764\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__41764\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__8496\ : InMux
    port map (
            O => \N__41761\,
            I => \N__41757\
        );

    \I__8495\ : InMux
    port map (
            O => \N__41760\,
            I => \N__41754\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__41757\,
            I => \N__41751\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__41754\,
            I => \N__41748\
        );

    \I__8492\ : Span4Mux_h
    port map (
            O => \N__41751\,
            I => \N__41745\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__41748\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__41745\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__8489\ : InMux
    port map (
            O => \N__41740\,
            I => \N__41736\
        );

    \I__8488\ : InMux
    port map (
            O => \N__41739\,
            I => \N__41733\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__41736\,
            I => \N__41730\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__41733\,
            I => \N__41727\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__41730\,
            I => \N__41724\
        );

    \I__8484\ : Odrv12
    port map (
            O => \N__41727\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__8483\ : Odrv4
    port map (
            O => \N__41724\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__41719\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__8481\ : InMux
    port map (
            O => \N__41716\,
            I => \N__41710\
        );

    \I__8480\ : InMux
    port map (
            O => \N__41715\,
            I => \N__41710\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__41710\,
            I => \N__41707\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__41707\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__8477\ : InMux
    port map (
            O => \N__41704\,
            I => \N__41700\
        );

    \I__8476\ : InMux
    port map (
            O => \N__41703\,
            I => \N__41697\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__41700\,
            I => \N__41692\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41692\
        );

    \I__8473\ : Odrv12
    port map (
            O => \N__41692\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__8472\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41683\
        );

    \I__8471\ : InMux
    port map (
            O => \N__41688\,
            I => \N__41683\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__41683\,
            I => \N__41680\
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__41680\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__41677\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__8467\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41671\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__41671\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__8465\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41665\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__41665\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__8463\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41658\
        );

    \I__8462\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41655\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41650\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__41655\,
            I => \N__41650\
        );

    \I__8459\ : Odrv12
    port map (
            O => \N__41650\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__8458\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41643\
        );

    \I__8457\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41640\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41635\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__41640\,
            I => \N__41635\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__41635\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__8453\ : CascadeMux
    port map (
            O => \N__41632\,
            I => \N__41629\
        );

    \I__8452\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41626\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__41626\,
            I => \N__41622\
        );

    \I__8450\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41619\
        );

    \I__8449\ : Span4Mux_h
    port map (
            O => \N__41622\,
            I => \N__41614\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__41619\,
            I => \N__41614\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__41614\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__8446\ : InMux
    port map (
            O => \N__41611\,
            I => \N__41608\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__41608\,
            I => \N__41604\
        );

    \I__8444\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41601\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__41604\,
            I => \N__41598\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__41601\,
            I => \N__41595\
        );

    \I__8441\ : Odrv4
    port map (
            O => \N__41598\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__8440\ : Odrv12
    port map (
            O => \N__41595\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__8439\ : InMux
    port map (
            O => \N__41590\,
            I => \N__41587\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__41587\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__8437\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41581\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__41581\,
            I => \N__41578\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__41578\,
            I => \N__41575\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__41575\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__8433\ : CascadeMux
    port map (
            O => \N__41572\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\
        );

    \I__8432\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41566\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__41566\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__8430\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41560\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__41560\,
            I => \N__41556\
        );

    \I__8428\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41553\
        );

    \I__8427\ : Span4Mux_h
    port map (
            O => \N__41556\,
            I => \N__41550\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__41553\,
            I => \N__41547\
        );

    \I__8425\ : Odrv4
    port map (
            O => \N__41550\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_15
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__41547\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_15
        );

    \I__8423\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41539\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__41539\,
            I => \N__41536\
        );

    \I__8421\ : Odrv4
    port map (
            O => \N__41536\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\
        );

    \I__8420\ : InMux
    port map (
            O => \N__41533\,
            I => \N__41530\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__41530\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__8418\ : InMux
    port map (
            O => \N__41527\,
            I => \N__41524\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__41524\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__8416\ : InMux
    port map (
            O => \N__41521\,
            I => \N__41518\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__41518\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__8414\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41512\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__41512\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__8412\ : InMux
    port map (
            O => \N__41509\,
            I => \N__41506\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__41506\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__8410\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41500\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__41500\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__8408\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41494\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__41494\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__8406\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41488\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__41488\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__8404\ : InMux
    port map (
            O => \N__41485\,
            I => \N__41482\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__41482\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__41479\,
            I => \N__41476\
        );

    \I__8401\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41473\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41470\
        );

    \I__8399\ : Span4Mux_v
    port map (
            O => \N__41470\,
            I => \N__41467\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__41467\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__8397\ : InMux
    port map (
            O => \N__41464\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__8396\ : InMux
    port map (
            O => \N__41461\,
            I => \N__41458\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__41458\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__8394\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41452\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__41452\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__8392\ : InMux
    port map (
            O => \N__41449\,
            I => \N__41446\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__41446\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__8390\ : InMux
    port map (
            O => \N__41443\,
            I => \N__41440\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__41440\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__8388\ : InMux
    port map (
            O => \N__41437\,
            I => \N__41434\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__41434\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__8386\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41428\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__41428\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__8384\ : InMux
    port map (
            O => \N__41425\,
            I => \N__41422\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__41422\,
            I => \N__41419\
        );

    \I__8382\ : Odrv12
    port map (
            O => \N__41419\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__8381\ : CascadeMux
    port map (
            O => \N__41416\,
            I => \N__41413\
        );

    \I__8380\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41410\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__41410\,
            I => \N__41407\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__41407\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__8377\ : InMux
    port map (
            O => \N__41404\,
            I => \N__41401\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__41401\,
            I => \N__41398\
        );

    \I__8375\ : Odrv4
    port map (
            O => \N__41398\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__8374\ : CascadeMux
    port map (
            O => \N__41395\,
            I => \N__41392\
        );

    \I__8373\ : InMux
    port map (
            O => \N__41392\,
            I => \N__41389\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__41389\,
            I => \N__41386\
        );

    \I__8371\ : Odrv4
    port map (
            O => \N__41386\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__8370\ : CascadeMux
    port map (
            O => \N__41383\,
            I => \N__41380\
        );

    \I__8369\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41377\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__41377\,
            I => \N__41374\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__41374\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8366\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41368\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__41368\,
            I => \N__41365\
        );

    \I__8364\ : Odrv12
    port map (
            O => \N__41365\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8363\ : CascadeMux
    port map (
            O => \N__41362\,
            I => \N__41359\
        );

    \I__8362\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41356\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__41356\,
            I => \N__41353\
        );

    \I__8360\ : Odrv4
    port map (
            O => \N__41353\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8359\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41347\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__41347\,
            I => \N__41344\
        );

    \I__8357\ : Odrv4
    port map (
            O => \N__41344\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__8356\ : CascadeMux
    port map (
            O => \N__41341\,
            I => \N__41338\
        );

    \I__8355\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41335\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__41335\,
            I => \N__41332\
        );

    \I__8353\ : Odrv4
    port map (
            O => \N__41332\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__41329\,
            I => \N__41326\
        );

    \I__8351\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41323\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41320\
        );

    \I__8349\ : Odrv4
    port map (
            O => \N__41320\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41314\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__41314\,
            I => \N__41311\
        );

    \I__8346\ : Odrv12
    port map (
            O => \N__41311\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__41308\,
            I => \N__41305\
        );

    \I__8344\ : InMux
    port map (
            O => \N__41305\,
            I => \N__41302\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__41302\,
            I => \N__41299\
        );

    \I__8342\ : Odrv12
    port map (
            O => \N__41299\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__8341\ : CascadeMux
    port map (
            O => \N__41296\,
            I => \N__41293\
        );

    \I__8340\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41290\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__41290\,
            I => \N__41287\
        );

    \I__8338\ : Odrv12
    port map (
            O => \N__41287\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__8337\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41281\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41278\
        );

    \I__8335\ : Odrv12
    port map (
            O => \N__41278\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__8334\ : InMux
    port map (
            O => \N__41275\,
            I => \N__41272\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__41272\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\
        );

    \I__8332\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41265\
        );

    \I__8331\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41262\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__41265\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__41262\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__8328\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41253\
        );

    \I__8327\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41250\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__41253\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__41250\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__8324\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41240\
        );

    \I__8323\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41237\
        );

    \I__8322\ : InMux
    port map (
            O => \N__41243\,
            I => \N__41234\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__41240\,
            I => \N__41231\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__41237\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__41234\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__8318\ : Odrv12
    port map (
            O => \N__41231\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__8317\ : InMux
    port map (
            O => \N__41224\,
            I => \N__41221\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__41221\,
            I => \N__41218\
        );

    \I__8315\ : Span4Mux_h
    port map (
            O => \N__41218\,
            I => \N__41214\
        );

    \I__8314\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41211\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__41214\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_21
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__41211\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_21
        );

    \I__8311\ : InMux
    port map (
            O => \N__41206\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\
        );

    \I__8310\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41200\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__41200\,
            I => \N__41197\
        );

    \I__8308\ : Span4Mux_h
    port map (
            O => \N__41197\,
            I => \N__41193\
        );

    \I__8307\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41190\
        );

    \I__8306\ : Odrv4
    port map (
            O => \N__41193\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_22
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__41190\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_22
        );

    \I__8304\ : InMux
    port map (
            O => \N__41185\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\
        );

    \I__8303\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41179\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__41179\,
            I => \N__41176\
        );

    \I__8301\ : Span4Mux_h
    port map (
            O => \N__41176\,
            I => \N__41172\
        );

    \I__8300\ : InMux
    port map (
            O => \N__41175\,
            I => \N__41169\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__41172\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_23
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__41169\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_23
        );

    \I__8297\ : InMux
    port map (
            O => \N__41164\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\
        );

    \I__8296\ : InMux
    port map (
            O => \N__41161\,
            I => \N__41158\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__41158\,
            I => \N__41154\
        );

    \I__8294\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41151\
        );

    \I__8293\ : Odrv12
    port map (
            O => \N__41154\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_24
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__41151\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_24
        );

    \I__8291\ : InMux
    port map (
            O => \N__41146\,
            I => \bfn_15_10_0_\
        );

    \I__8290\ : InMux
    port map (
            O => \N__41143\,
            I => \N__41140\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__41140\,
            I => \N__41137\
        );

    \I__8288\ : Span12Mux_s9_v
    port map (
            O => \N__41137\,
            I => \N__41133\
        );

    \I__8287\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41130\
        );

    \I__8286\ : Odrv12
    port map (
            O => \N__41133\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_25
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__41130\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_25
        );

    \I__8284\ : InMux
    port map (
            O => \N__41125\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\
        );

    \I__8283\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41119\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__41119\,
            I => \N__41115\
        );

    \I__8281\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41112\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__41115\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_26
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__41112\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_26
        );

    \I__8278\ : InMux
    port map (
            O => \N__41107\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\
        );

    \I__8277\ : InMux
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__41101\,
            I => \N__41097\
        );

    \I__8275\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41094\
        );

    \I__8274\ : Odrv4
    port map (
            O => \N__41097\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_27
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__41094\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_27
        );

    \I__8272\ : InMux
    port map (
            O => \N__41089\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\
        );

    \I__8271\ : InMux
    port map (
            O => \N__41086\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\
        );

    \I__8270\ : InMux
    port map (
            O => \N__41083\,
            I => \N__41080\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__41080\,
            I => \N__41076\
        );

    \I__8268\ : InMux
    port map (
            O => \N__41079\,
            I => \N__41073\
        );

    \I__8267\ : Span4Mux_h
    port map (
            O => \N__41076\,
            I => \N__41070\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__41073\,
            I => \N__41067\
        );

    \I__8265\ : Odrv4
    port map (
            O => \N__41070\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_13
        );

    \I__8264\ : Odrv4
    port map (
            O => \N__41067\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_13
        );

    \I__8263\ : InMux
    port map (
            O => \N__41062\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\
        );

    \I__8262\ : InMux
    port map (
            O => \N__41059\,
            I => \N__41056\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41052\
        );

    \I__8260\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41049\
        );

    \I__8259\ : Span4Mux_h
    port map (
            O => \N__41052\,
            I => \N__41046\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__41049\,
            I => \N__41043\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__41046\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_14
        );

    \I__8256\ : Odrv4
    port map (
            O => \N__41043\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_14
        );

    \I__8255\ : InMux
    port map (
            O => \N__41038\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\
        );

    \I__8254\ : InMux
    port map (
            O => \N__41035\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\
        );

    \I__8253\ : InMux
    port map (
            O => \N__41032\,
            I => \N__41028\
        );

    \I__8252\ : InMux
    port map (
            O => \N__41031\,
            I => \N__41025\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41022\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__41019\
        );

    \I__8249\ : Span4Mux_h
    port map (
            O => \N__41022\,
            I => \N__41016\
        );

    \I__8248\ : Span4Mux_h
    port map (
            O => \N__41019\,
            I => \N__41013\
        );

    \I__8247\ : Odrv4
    port map (
            O => \N__41016\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_16
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__41013\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_16
        );

    \I__8245\ : InMux
    port map (
            O => \N__41008\,
            I => \bfn_15_9_0_\
        );

    \I__8244\ : InMux
    port map (
            O => \N__41005\,
            I => \N__41001\
        );

    \I__8243\ : InMux
    port map (
            O => \N__41004\,
            I => \N__40998\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__41001\,
            I => \N__40995\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__40998\,
            I => \N__40992\
        );

    \I__8240\ : Span4Mux_h
    port map (
            O => \N__40995\,
            I => \N__40989\
        );

    \I__8239\ : Span4Mux_h
    port map (
            O => \N__40992\,
            I => \N__40986\
        );

    \I__8238\ : Odrv4
    port map (
            O => \N__40989\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_17
        );

    \I__8237\ : Odrv4
    port map (
            O => \N__40986\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_17
        );

    \I__8236\ : InMux
    port map (
            O => \N__40981\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\
        );

    \I__8235\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40974\
        );

    \I__8234\ : InMux
    port map (
            O => \N__40977\,
            I => \N__40971\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40966\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__40971\,
            I => \N__40966\
        );

    \I__8231\ : Span4Mux_h
    port map (
            O => \N__40966\,
            I => \N__40963\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__40963\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_18
        );

    \I__8229\ : InMux
    port map (
            O => \N__40960\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\
        );

    \I__8228\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40953\
        );

    \I__8227\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40950\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__40953\,
            I => \N__40947\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__40950\,
            I => \N__40944\
        );

    \I__8224\ : Span4Mux_h
    port map (
            O => \N__40947\,
            I => \N__40941\
        );

    \I__8223\ : Span4Mux_v
    port map (
            O => \N__40944\,
            I => \N__40938\
        );

    \I__8222\ : Odrv4
    port map (
            O => \N__40941\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_19
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__40938\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_19
        );

    \I__8220\ : InMux
    port map (
            O => \N__40933\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\
        );

    \I__8219\ : InMux
    port map (
            O => \N__40930\,
            I => \N__40927\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__40927\,
            I => \N__40924\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__40924\,
            I => \N__40920\
        );

    \I__8216\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40917\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__40920\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_20
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__40917\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_20
        );

    \I__8213\ : InMux
    port map (
            O => \N__40912\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\
        );

    \I__8212\ : InMux
    port map (
            O => \N__40909\,
            I => \N__40906\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__40906\,
            I => \N__40902\
        );

    \I__8210\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40899\
        );

    \I__8209\ : Span4Mux_h
    port map (
            O => \N__40902\,
            I => \N__40896\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__40899\,
            I => \N__40893\
        );

    \I__8207\ : Odrv4
    port map (
            O => \N__40896\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_4
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__40893\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_4
        );

    \I__8205\ : InMux
    port map (
            O => \N__40888\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\
        );

    \I__8204\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40882\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__40882\,
            I => \N__40878\
        );

    \I__8202\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40875\
        );

    \I__8201\ : Span4Mux_h
    port map (
            O => \N__40878\,
            I => \N__40872\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__40875\,
            I => \N__40869\
        );

    \I__8199\ : Odrv4
    port map (
            O => \N__40872\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_5
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__40869\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_5
        );

    \I__8197\ : InMux
    port map (
            O => \N__40864\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\
        );

    \I__8196\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40858\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__40858\,
            I => \N__40854\
        );

    \I__8194\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40851\
        );

    \I__8193\ : Span4Mux_h
    port map (
            O => \N__40854\,
            I => \N__40848\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__40851\,
            I => \N__40845\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__40848\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_6
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__40845\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_6
        );

    \I__8189\ : InMux
    port map (
            O => \N__40840\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\
        );

    \I__8188\ : InMux
    port map (
            O => \N__40837\,
            I => \N__40834\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__40834\,
            I => \N__40830\
        );

    \I__8186\ : InMux
    port map (
            O => \N__40833\,
            I => \N__40827\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__40830\,
            I => \N__40824\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__40827\,
            I => \N__40821\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__40824\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_7
        );

    \I__8182\ : Odrv4
    port map (
            O => \N__40821\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_7
        );

    \I__8181\ : InMux
    port map (
            O => \N__40816\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\
        );

    \I__8180\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40809\
        );

    \I__8179\ : InMux
    port map (
            O => \N__40812\,
            I => \N__40806\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__40809\,
            I => \N__40803\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__40806\,
            I => \N__40798\
        );

    \I__8176\ : Span4Mux_h
    port map (
            O => \N__40803\,
            I => \N__40798\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__40798\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_8
        );

    \I__8174\ : InMux
    port map (
            O => \N__40795\,
            I => \bfn_15_8_0_\
        );

    \I__8173\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40789\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__40789\,
            I => \N__40785\
        );

    \I__8171\ : InMux
    port map (
            O => \N__40788\,
            I => \N__40782\
        );

    \I__8170\ : Span4Mux_h
    port map (
            O => \N__40785\,
            I => \N__40779\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__40782\,
            I => \N__40776\
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__40779\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_9
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__40776\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_9
        );

    \I__8166\ : InMux
    port map (
            O => \N__40771\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\
        );

    \I__8165\ : InMux
    port map (
            O => \N__40768\,
            I => \N__40765\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__40765\,
            I => \N__40761\
        );

    \I__8163\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40758\
        );

    \I__8162\ : Span4Mux_v
    port map (
            O => \N__40761\,
            I => \N__40755\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__40758\,
            I => \N__40752\
        );

    \I__8160\ : Odrv4
    port map (
            O => \N__40755\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_10
        );

    \I__8159\ : Odrv4
    port map (
            O => \N__40752\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_10
        );

    \I__8158\ : InMux
    port map (
            O => \N__40747\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\
        );

    \I__8157\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40741\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40737\
        );

    \I__8155\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40734\
        );

    \I__8154\ : Span4Mux_v
    port map (
            O => \N__40737\,
            I => \N__40731\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__40734\,
            I => \N__40728\
        );

    \I__8152\ : Odrv4
    port map (
            O => \N__40731\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_11
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__40728\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_11
        );

    \I__8150\ : InMux
    port map (
            O => \N__40723\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\
        );

    \I__8149\ : InMux
    port map (
            O => \N__40720\,
            I => \N__40717\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__40717\,
            I => \N__40713\
        );

    \I__8147\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40710\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__40713\,
            I => \N__40707\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__40710\,
            I => \N__40704\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__40707\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_12
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__40704\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_12
        );

    \I__8142\ : InMux
    port map (
            O => \N__40699\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\
        );

    \I__8141\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40693\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__40693\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\
        );

    \I__8139\ : CascadeMux
    port map (
            O => \N__40690\,
            I => \N__40687\
        );

    \I__8138\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40684\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__40684\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\
        );

    \I__8136\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40678\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__40678\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\
        );

    \I__8134\ : InMux
    port map (
            O => \N__40675\,
            I => \N__40672\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__40672\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\
        );

    \I__8132\ : InMux
    port map (
            O => \N__40669\,
            I => \N__40666\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__40666\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\
        );

    \I__8130\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40660\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__40660\,
            I => \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\
        );

    \I__8128\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40654\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__40654\,
            I => \N__40650\
        );

    \I__8126\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40647\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__40650\,
            I => \N__40644\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__40647\,
            I => \N__40641\
        );

    \I__8123\ : Odrv4
    port map (
            O => \N__40644\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_1
        );

    \I__8122\ : Odrv4
    port map (
            O => \N__40641\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_1
        );

    \I__8121\ : InMux
    port map (
            O => \N__40636\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\
        );

    \I__8120\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40630\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__40630\,
            I => \N__40626\
        );

    \I__8118\ : InMux
    port map (
            O => \N__40629\,
            I => \N__40623\
        );

    \I__8117\ : Span4Mux_v
    port map (
            O => \N__40626\,
            I => \N__40620\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__40623\,
            I => \N__40617\
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__40620\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_2
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__40617\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_2
        );

    \I__8113\ : InMux
    port map (
            O => \N__40612\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\
        );

    \I__8112\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40606\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__40606\,
            I => \N__40602\
        );

    \I__8110\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40599\
        );

    \I__8109\ : Span4Mux_v
    port map (
            O => \N__40602\,
            I => \N__40596\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__40599\,
            I => \N__40593\
        );

    \I__8107\ : Odrv4
    port map (
            O => \N__40596\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_3
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__40593\,
            I => phase_controller_inst1_stoper_hc_target_ticks_1_i_3
        );

    \I__8105\ : InMux
    port map (
            O => \N__40588\,
            I => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__40585\,
            I => \N__40582\
        );

    \I__8103\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40579\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__40579\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\
        );

    \I__8101\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__40573\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\
        );

    \I__8099\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40567\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__40567\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__40564\,
            I => \N__40561\
        );

    \I__8096\ : InMux
    port map (
            O => \N__40561\,
            I => \N__40558\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__40558\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\
        );

    \I__8094\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40552\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__40552\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\
        );

    \I__8092\ : InMux
    port map (
            O => \N__40549\,
            I => \N__40546\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__40546\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\
        );

    \I__8090\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40540\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__40540\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\
        );

    \I__8088\ : InMux
    port map (
            O => \N__40537\,
            I => \N__40534\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__40534\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\
        );

    \I__8086\ : InMux
    port map (
            O => \N__40531\,
            I => \N__40528\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__40528\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\
        );

    \I__8084\ : CascadeMux
    port map (
            O => \N__40525\,
            I => \current_shift_inst.control_input_31_cascade_\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__40522\,
            I => \N__40519\
        );

    \I__8082\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40516\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__40516\,
            I => \N__40513\
        );

    \I__8080\ : Odrv4
    port map (
            O => \N__40513\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__8079\ : CascadeMux
    port map (
            O => \N__40510\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\
        );

    \I__8078\ : InMux
    port map (
            O => \N__40507\,
            I => \N__40504\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__40504\,
            I => \N__40500\
        );

    \I__8076\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40497\
        );

    \I__8075\ : Span4Mux_h
    port map (
            O => \N__40500\,
            I => \N__40494\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__40497\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__40494\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__8072\ : CascadeMux
    port map (
            O => \N__40489\,
            I => \N__40486\
        );

    \I__8071\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40483\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__40483\,
            I => \N__40479\
        );

    \I__8069\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40476\
        );

    \I__8068\ : Span4Mux_h
    port map (
            O => \N__40479\,
            I => \N__40473\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__40476\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__8066\ : Odrv4
    port map (
            O => \N__40473\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__40468\,
            I => \N__40464\
        );

    \I__8064\ : InMux
    port map (
            O => \N__40467\,
            I => \N__40461\
        );

    \I__8063\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40458\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__40461\,
            I => \N__40455\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__40458\,
            I => \N__40450\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__40455\,
            I => \N__40450\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__40450\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__40447\,
            I => \N__40444\
        );

    \I__8057\ : InMux
    port map (
            O => \N__40444\,
            I => \N__40441\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__40441\,
            I => \N__40437\
        );

    \I__8055\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40434\
        );

    \I__8054\ : Span4Mux_h
    port map (
            O => \N__40437\,
            I => \N__40431\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__40434\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__40431\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__8051\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40423\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__40423\,
            I => \N__40419\
        );

    \I__8049\ : InMux
    port map (
            O => \N__40422\,
            I => \N__40416\
        );

    \I__8048\ : Span4Mux_v
    port map (
            O => \N__40419\,
            I => \N__40411\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__40416\,
            I => \N__40411\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__40411\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__8045\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40402\
        );

    \I__8044\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40402\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__40402\,
            I => \N__40399\
        );

    \I__8042\ : Odrv4
    port map (
            O => \N__40399\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__40396\,
            I => \N__40393\
        );

    \I__8040\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40387\
        );

    \I__8039\ : InMux
    port map (
            O => \N__40392\,
            I => \N__40387\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__40387\,
            I => \N__40384\
        );

    \I__8037\ : Span4Mux_h
    port map (
            O => \N__40384\,
            I => \N__40381\
        );

    \I__8036\ : Odrv4
    port map (
            O => \N__40381\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__8035\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40372\
        );

    \I__8034\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40372\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__40372\,
            I => \N__40369\
        );

    \I__8032\ : Odrv12
    port map (
            O => \N__40369\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__8031\ : ClkMux
    port map (
            O => \N__40366\,
            I => \N__40363\
        );

    \I__8030\ : GlobalMux
    port map (
            O => \N__40363\,
            I => \N__40360\
        );

    \I__8029\ : gio2CtrlBuf
    port map (
            O => \N__40360\,
            I => delay_hc_input_c_g
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__40357\,
            I => \N__40354\
        );

    \I__8027\ : InMux
    port map (
            O => \N__40354\,
            I => \N__40351\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__40351\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\
        );

    \I__8025\ : InMux
    port map (
            O => \N__40348\,
            I => \N__40345\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__40345\,
            I => \N__40342\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__40342\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__8022\ : InMux
    port map (
            O => \N__40339\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__8021\ : InMux
    port map (
            O => \N__40336\,
            I => \N__40333\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__40333\,
            I => \N__40330\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__40330\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__8018\ : InMux
    port map (
            O => \N__40327\,
            I => \bfn_14_22_0_\
        );

    \I__8017\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40321\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40318\
        );

    \I__8015\ : Odrv4
    port map (
            O => \N__40318\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__8014\ : InMux
    port map (
            O => \N__40315\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__8013\ : InMux
    port map (
            O => \N__40312\,
            I => \N__40309\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__40309\,
            I => \N__40306\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__40306\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__8010\ : InMux
    port map (
            O => \N__40303\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__8009\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40297\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__40297\,
            I => \N__40294\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__40294\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__8006\ : InMux
    port map (
            O => \N__40291\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__8005\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40285\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__40285\,
            I => \N__40282\
        );

    \I__8003\ : Odrv4
    port map (
            O => \N__40282\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__8002\ : InMux
    port map (
            O => \N__40279\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__8001\ : InMux
    port map (
            O => \N__40276\,
            I => \N__40273\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__40273\,
            I => \N__40270\
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__40270\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__7998\ : InMux
    port map (
            O => \N__40267\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__7997\ : InMux
    port map (
            O => \N__40264\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__7996\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40258\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__40258\,
            I => \N__40255\
        );

    \I__7994\ : Odrv4
    port map (
            O => \N__40255\,
            I => \current_shift_inst.control_input_31\
        );

    \I__7993\ : InMux
    port map (
            O => \N__40252\,
            I => \N__40249\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__40249\,
            I => \N__40246\
        );

    \I__7991\ : Odrv4
    port map (
            O => \N__40246\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__7990\ : InMux
    port map (
            O => \N__40243\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__7989\ : InMux
    port map (
            O => \N__40240\,
            I => \N__40237\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__40237\,
            I => \N__40234\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__40234\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__7986\ : InMux
    port map (
            O => \N__40231\,
            I => \bfn_14_21_0_\
        );

    \I__7985\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40225\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__40225\,
            I => \N__40222\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__40222\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__7982\ : InMux
    port map (
            O => \N__40219\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__7981\ : InMux
    port map (
            O => \N__40216\,
            I => \N__40213\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__7979\ : Odrv4
    port map (
            O => \N__40210\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__7978\ : InMux
    port map (
            O => \N__40207\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__7977\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40201\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__40201\,
            I => \N__40198\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__40198\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__7974\ : InMux
    port map (
            O => \N__40195\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__7973\ : InMux
    port map (
            O => \N__40192\,
            I => \N__40189\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__40189\,
            I => \N__40186\
        );

    \I__7971\ : Odrv4
    port map (
            O => \N__40186\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__7970\ : InMux
    port map (
            O => \N__40183\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__7969\ : InMux
    port map (
            O => \N__40180\,
            I => \N__40177\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__40177\,
            I => \N__40174\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__40174\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__7966\ : InMux
    port map (
            O => \N__40171\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__7965\ : CascadeMux
    port map (
            O => \N__40168\,
            I => \N__40165\
        );

    \I__7964\ : InMux
    port map (
            O => \N__40165\,
            I => \N__40162\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__40162\,
            I => \N__40159\
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__40159\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__7961\ : InMux
    port map (
            O => \N__40156\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__40153\,
            I => \N__40150\
        );

    \I__7959\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40147\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__40147\,
            I => \N__40144\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__40144\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__7956\ : InMux
    port map (
            O => \N__40141\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__7955\ : InMux
    port map (
            O => \N__40138\,
            I => \N__40135\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__40132\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__7952\ : InMux
    port map (
            O => \N__40129\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__7951\ : InMux
    port map (
            O => \N__40126\,
            I => \N__40123\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__40123\,
            I => \N__40120\
        );

    \I__7949\ : Odrv4
    port map (
            O => \N__40120\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__7948\ : InMux
    port map (
            O => \N__40117\,
            I => \bfn_14_20_0_\
        );

    \I__7947\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40111\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__40111\,
            I => \N__40108\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__40108\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__7944\ : InMux
    port map (
            O => \N__40105\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__7943\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40099\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__40099\,
            I => \N__40096\
        );

    \I__7941\ : Odrv4
    port map (
            O => \N__40096\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__7940\ : InMux
    port map (
            O => \N__40093\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__7939\ : InMux
    port map (
            O => \N__40090\,
            I => \N__40087\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__40087\,
            I => \N__40084\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__40084\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__7936\ : InMux
    port map (
            O => \N__40081\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__7935\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40075\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__40075\,
            I => \N__40072\
        );

    \I__7933\ : Odrv4
    port map (
            O => \N__40072\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__7932\ : InMux
    port map (
            O => \N__40069\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__7931\ : InMux
    port map (
            O => \N__40066\,
            I => \N__40063\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__40063\,
            I => \N__40060\
        );

    \I__7929\ : Odrv4
    port map (
            O => \N__40060\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__7928\ : InMux
    port map (
            O => \N__40057\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__40054\,
            I => \N__40051\
        );

    \I__7926\ : InMux
    port map (
            O => \N__40051\,
            I => \N__40048\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__40048\,
            I => \N__40045\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__40045\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__7923\ : InMux
    port map (
            O => \N__40042\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__7922\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40036\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__40036\,
            I => \N__40033\
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__40033\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7919\ : InMux
    port map (
            O => \N__40030\,
            I => \N__40027\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__40027\,
            I => \N__40024\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__40024\,
            I => \current_shift_inst.control_input_1\
        );

    \I__7916\ : InMux
    port map (
            O => \N__40021\,
            I => \N__40018\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__40018\,
            I => \N__40015\
        );

    \I__7914\ : Odrv4
    port map (
            O => \N__40015\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__7913\ : InMux
    port map (
            O => \N__40012\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__7912\ : InMux
    port map (
            O => \N__40009\,
            I => \N__40006\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__40006\,
            I => \N__40003\
        );

    \I__7910\ : Odrv4
    port map (
            O => \N__40003\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__7909\ : InMux
    port map (
            O => \N__40000\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__7908\ : InMux
    port map (
            O => \N__39997\,
            I => \N__39994\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__39994\,
            I => \N__39991\
        );

    \I__7906\ : Odrv4
    port map (
            O => \N__39991\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__7905\ : InMux
    port map (
            O => \N__39988\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__7904\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39982\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__39982\,
            I => \N__39979\
        );

    \I__7902\ : Span4Mux_h
    port map (
            O => \N__39979\,
            I => \N__39976\
        );

    \I__7901\ : Odrv4
    port map (
            O => \N__39976\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__7900\ : InMux
    port map (
            O => \N__39973\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__7899\ : InMux
    port map (
            O => \N__39970\,
            I => \N__39967\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__39967\,
            I => \N__39964\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__39964\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__7896\ : InMux
    port map (
            O => \N__39961\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__7895\ : CascadeMux
    port map (
            O => \N__39958\,
            I => \N__39954\
        );

    \I__7894\ : CascadeMux
    port map (
            O => \N__39957\,
            I => \N__39951\
        );

    \I__7893\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39945\
        );

    \I__7892\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39945\
        );

    \I__7891\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39942\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__39945\,
            I => \N__39939\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__39942\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__7888\ : Odrv12
    port map (
            O => \N__39939\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__7887\ : InMux
    port map (
            O => \N__39934\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__7886\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39925\
        );

    \I__7885\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39925\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__39925\,
            I => \N__39921\
        );

    \I__7883\ : InMux
    port map (
            O => \N__39924\,
            I => \N__39918\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__39921\,
            I => \N__39915\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__39918\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__39915\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__7879\ : InMux
    port map (
            O => \N__39910\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__7878\ : CascadeMux
    port map (
            O => \N__39907\,
            I => \N__39904\
        );

    \I__7877\ : InMux
    port map (
            O => \N__39904\,
            I => \N__39900\
        );

    \I__7876\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39897\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__39900\,
            I => \N__39891\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__39897\,
            I => \N__39891\
        );

    \I__7873\ : InMux
    port map (
            O => \N__39896\,
            I => \N__39888\
        );

    \I__7872\ : Span4Mux_v
    port map (
            O => \N__39891\,
            I => \N__39885\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__39888\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__39885\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__7869\ : InMux
    port map (
            O => \N__39880\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__7868\ : CascadeMux
    port map (
            O => \N__39877\,
            I => \N__39873\
        );

    \I__7867\ : CascadeMux
    port map (
            O => \N__39876\,
            I => \N__39870\
        );

    \I__7866\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39866\
        );

    \I__7865\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39863\
        );

    \I__7864\ : InMux
    port map (
            O => \N__39869\,
            I => \N__39860\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__39866\,
            I => \N__39855\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__39863\,
            I => \N__39855\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__39860\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7860\ : Odrv12
    port map (
            O => \N__39855\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7859\ : InMux
    port map (
            O => \N__39850\,
            I => \bfn_14_18_0_\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__39847\,
            I => \N__39844\
        );

    \I__7857\ : InMux
    port map (
            O => \N__39844\,
            I => \N__39841\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__39841\,
            I => \N__39836\
        );

    \I__7855\ : InMux
    port map (
            O => \N__39840\,
            I => \N__39833\
        );

    \I__7854\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39830\
        );

    \I__7853\ : Sp12to4
    port map (
            O => \N__39836\,
            I => \N__39825\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__39833\,
            I => \N__39825\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__39830\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7850\ : Odrv12
    port map (
            O => \N__39825\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7849\ : InMux
    port map (
            O => \N__39820\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__7848\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39813\
        );

    \I__7847\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39810\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__39813\,
            I => \N__39807\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__39810\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7844\ : Odrv12
    port map (
            O => \N__39807\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__39802\,
            I => \N__39799\
        );

    \I__7842\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39794\
        );

    \I__7841\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39791\
        );

    \I__7840\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39788\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39783\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__39791\,
            I => \N__39783\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__39788\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7836\ : Odrv12
    port map (
            O => \N__39783\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7835\ : InMux
    port map (
            O => \N__39778\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__7834\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39772\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__39772\,
            I => \N__39768\
        );

    \I__7832\ : InMux
    port map (
            O => \N__39771\,
            I => \N__39765\
        );

    \I__7831\ : Span4Mux_v
    port map (
            O => \N__39768\,
            I => \N__39762\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__39765\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__39762\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__39757\,
            I => \N__39754\
        );

    \I__7827\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39749\
        );

    \I__7826\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39746\
        );

    \I__7825\ : InMux
    port map (
            O => \N__39752\,
            I => \N__39743\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__39749\,
            I => \N__39738\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__39746\,
            I => \N__39738\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__39743\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7821\ : Odrv12
    port map (
            O => \N__39738\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7820\ : InMux
    port map (
            O => \N__39733\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__7819\ : InMux
    port map (
            O => \N__39730\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__7818\ : CascadeMux
    port map (
            O => \N__39727\,
            I => \N__39723\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__39726\,
            I => \N__39720\
        );

    \I__7816\ : InMux
    port map (
            O => \N__39723\,
            I => \N__39714\
        );

    \I__7815\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39714\
        );

    \I__7814\ : InMux
    port map (
            O => \N__39719\,
            I => \N__39711\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__39714\,
            I => \N__39708\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__39711\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__7811\ : Odrv12
    port map (
            O => \N__39708\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__7810\ : InMux
    port map (
            O => \N__39703\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__39700\,
            I => \N__39696\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__39699\,
            I => \N__39693\
        );

    \I__7807\ : InMux
    port map (
            O => \N__39696\,
            I => \N__39688\
        );

    \I__7806\ : InMux
    port map (
            O => \N__39693\,
            I => \N__39688\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__39688\,
            I => \N__39684\
        );

    \I__7804\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39681\
        );

    \I__7803\ : Span4Mux_v
    port map (
            O => \N__39684\,
            I => \N__39678\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__39681\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__7801\ : Odrv4
    port map (
            O => \N__39678\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__7800\ : InMux
    port map (
            O => \N__39673\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__39670\,
            I => \N__39667\
        );

    \I__7798\ : InMux
    port map (
            O => \N__39667\,
            I => \N__39662\
        );

    \I__7797\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39659\
        );

    \I__7796\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39656\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__39662\,
            I => \N__39651\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__39659\,
            I => \N__39651\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__39656\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__7792\ : Odrv12
    port map (
            O => \N__39651\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__7791\ : InMux
    port map (
            O => \N__39646\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__39643\,
            I => \N__39640\
        );

    \I__7789\ : InMux
    port map (
            O => \N__39640\,
            I => \N__39637\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__39637\,
            I => \N__39632\
        );

    \I__7787\ : InMux
    port map (
            O => \N__39636\,
            I => \N__39629\
        );

    \I__7786\ : InMux
    port map (
            O => \N__39635\,
            I => \N__39626\
        );

    \I__7785\ : Sp12to4
    port map (
            O => \N__39632\,
            I => \N__39621\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__39629\,
            I => \N__39621\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__39626\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7782\ : Odrv12
    port map (
            O => \N__39621\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7781\ : InMux
    port map (
            O => \N__39616\,
            I => \bfn_14_17_0_\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__39613\,
            I => \N__39610\
        );

    \I__7779\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39607\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__39607\,
            I => \N__39602\
        );

    \I__7777\ : InMux
    port map (
            O => \N__39606\,
            I => \N__39599\
        );

    \I__7776\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39596\
        );

    \I__7775\ : Sp12to4
    port map (
            O => \N__39602\,
            I => \N__39591\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__39599\,
            I => \N__39591\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__39596\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7772\ : Odrv12
    port map (
            O => \N__39591\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7771\ : InMux
    port map (
            O => \N__39586\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__7770\ : InMux
    port map (
            O => \N__39583\,
            I => \N__39576\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39582\,
            I => \N__39576\
        );

    \I__7768\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39573\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__39576\,
            I => \N__39570\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__39573\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__7765\ : Odrv12
    port map (
            O => \N__39570\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__7764\ : InMux
    port map (
            O => \N__39565\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__7763\ : InMux
    port map (
            O => \N__39562\,
            I => \N__39555\
        );

    \I__7762\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39555\
        );

    \I__7761\ : InMux
    port map (
            O => \N__39560\,
            I => \N__39552\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__39555\,
            I => \N__39549\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__39552\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__7758\ : Odrv12
    port map (
            O => \N__39549\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__7757\ : InMux
    port map (
            O => \N__39544\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__39541\,
            I => \N__39537\
        );

    \I__7755\ : CascadeMux
    port map (
            O => \N__39540\,
            I => \N__39534\
        );

    \I__7754\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39528\
        );

    \I__7753\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39528\
        );

    \I__7752\ : InMux
    port map (
            O => \N__39533\,
            I => \N__39525\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__39528\,
            I => \N__39522\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__39525\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__7749\ : Odrv12
    port map (
            O => \N__39522\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__7748\ : InMux
    port map (
            O => \N__39517\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__7747\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39508\
        );

    \I__7746\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39508\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__39508\,
            I => \N__39504\
        );

    \I__7744\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39501\
        );

    \I__7743\ : Span4Mux_v
    port map (
            O => \N__39504\,
            I => \N__39498\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__39501\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__7741\ : Odrv4
    port map (
            O => \N__39498\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__7740\ : InMux
    port map (
            O => \N__39493\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__39490\,
            I => \N__39486\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__39489\,
            I => \N__39483\
        );

    \I__7737\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39477\
        );

    \I__7736\ : InMux
    port map (
            O => \N__39483\,
            I => \N__39477\
        );

    \I__7735\ : InMux
    port map (
            O => \N__39482\,
            I => \N__39474\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__39477\,
            I => \N__39471\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__39474\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__7732\ : Odrv12
    port map (
            O => \N__39471\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__7731\ : InMux
    port map (
            O => \N__39466\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__39463\,
            I => \N__39459\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__39462\,
            I => \N__39456\
        );

    \I__7728\ : InMux
    port map (
            O => \N__39459\,
            I => \N__39451\
        );

    \I__7727\ : InMux
    port map (
            O => \N__39456\,
            I => \N__39451\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__39451\,
            I => \N__39447\
        );

    \I__7725\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39444\
        );

    \I__7724\ : Span4Mux_v
    port map (
            O => \N__39447\,
            I => \N__39441\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__39444\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__39441\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__7721\ : InMux
    port map (
            O => \N__39436\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__7720\ : CascadeMux
    port map (
            O => \N__39433\,
            I => \N__39430\
        );

    \I__7719\ : InMux
    port map (
            O => \N__39430\,
            I => \N__39426\
        );

    \I__7718\ : InMux
    port map (
            O => \N__39429\,
            I => \N__39423\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__39426\,
            I => \N__39417\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__39423\,
            I => \N__39417\
        );

    \I__7715\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39414\
        );

    \I__7714\ : Span4Mux_v
    port map (
            O => \N__39417\,
            I => \N__39411\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__39414\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__7712\ : Odrv4
    port map (
            O => \N__39411\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__7711\ : InMux
    port map (
            O => \N__39406\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__39403\,
            I => \N__39400\
        );

    \I__7709\ : InMux
    port map (
            O => \N__39400\,
            I => \N__39395\
        );

    \I__7708\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39392\
        );

    \I__7707\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39389\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__39395\,
            I => \N__39384\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__39392\,
            I => \N__39384\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__39389\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7703\ : Odrv12
    port map (
            O => \N__39384\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7702\ : InMux
    port map (
            O => \N__39379\,
            I => \bfn_14_16_0_\
        );

    \I__7701\ : CascadeMux
    port map (
            O => \N__39376\,
            I => \N__39373\
        );

    \I__7700\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39370\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__39370\,
            I => \N__39365\
        );

    \I__7698\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39362\
        );

    \I__7697\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39359\
        );

    \I__7696\ : Sp12to4
    port map (
            O => \N__39365\,
            I => \N__39354\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__39362\,
            I => \N__39354\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__39359\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7693\ : Odrv12
    port map (
            O => \N__39354\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7692\ : InMux
    port map (
            O => \N__39349\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__39346\,
            I => \N__39343\
        );

    \I__7690\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39339\
        );

    \I__7689\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39336\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__39339\,
            I => \N__39330\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__39336\,
            I => \N__39330\
        );

    \I__7686\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39327\
        );

    \I__7685\ : Span4Mux_v
    port map (
            O => \N__39330\,
            I => \N__39324\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__39327\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__39324\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__7682\ : InMux
    port map (
            O => \N__39319\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__7681\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39310\
        );

    \I__7680\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39310\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__39310\,
            I => \N__39306\
        );

    \I__7678\ : InMux
    port map (
            O => \N__39309\,
            I => \N__39303\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__39306\,
            I => \N__39300\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__39303\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__39300\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__7674\ : InMux
    port map (
            O => \N__39295\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__7673\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39286\
        );

    \I__7672\ : InMux
    port map (
            O => \N__39291\,
            I => \N__39286\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39282\
        );

    \I__7670\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39279\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__39282\,
            I => \N__39276\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__39279\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__39276\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__7666\ : InMux
    port map (
            O => \N__39271\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__7665\ : InMux
    port map (
            O => \N__39268\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__7664\ : InMux
    port map (
            O => \N__39265\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__7663\ : InMux
    port map (
            O => \N__39262\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__7662\ : InMux
    port map (
            O => \N__39259\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__7661\ : InMux
    port map (
            O => \N__39256\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__7660\ : InMux
    port map (
            O => \N__39253\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__7659\ : CascadeMux
    port map (
            O => \N__39250\,
            I => \N__39246\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__39249\,
            I => \N__39243\
        );

    \I__7657\ : InMux
    port map (
            O => \N__39246\,
            I => \N__39238\
        );

    \I__7656\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39238\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__39238\,
            I => \N__39234\
        );

    \I__7654\ : InMux
    port map (
            O => \N__39237\,
            I => \N__39231\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__39234\,
            I => \N__39228\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__39231\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7651\ : Odrv4
    port map (
            O => \N__39228\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7650\ : InMux
    port map (
            O => \N__39223\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__7649\ : CascadeMux
    port map (
            O => \N__39220\,
            I => \N__39216\
        );

    \I__7648\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39213\
        );

    \I__7647\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39210\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__39213\,
            I => \N__39204\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__39210\,
            I => \N__39204\
        );

    \I__7644\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39201\
        );

    \I__7643\ : Span4Mux_v
    port map (
            O => \N__39204\,
            I => \N__39198\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__39201\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7641\ : Odrv4
    port map (
            O => \N__39198\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7640\ : InMux
    port map (
            O => \N__39193\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__7639\ : InMux
    port map (
            O => \N__39190\,
            I => \bfn_14_13_0_\
        );

    \I__7638\ : InMux
    port map (
            O => \N__39187\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__7637\ : InMux
    port map (
            O => \N__39184\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__7636\ : InMux
    port map (
            O => \N__39181\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__7635\ : InMux
    port map (
            O => \N__39178\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__7634\ : InMux
    port map (
            O => \N__39175\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__7633\ : InMux
    port map (
            O => \N__39172\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__7632\ : InMux
    port map (
            O => \N__39169\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__7631\ : InMux
    port map (
            O => \N__39166\,
            I => \bfn_14_14_0_\
        );

    \I__7630\ : InMux
    port map (
            O => \N__39163\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__7629\ : InMux
    port map (
            O => \N__39160\,
            I => \bfn_14_12_0_\
        );

    \I__7628\ : InMux
    port map (
            O => \N__39157\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__7627\ : InMux
    port map (
            O => \N__39154\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__7626\ : InMux
    port map (
            O => \N__39151\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__7625\ : InMux
    port map (
            O => \N__39148\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__7624\ : InMux
    port map (
            O => \N__39145\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__7623\ : InMux
    port map (
            O => \N__39142\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__7622\ : InMux
    port map (
            O => \N__39139\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__7621\ : InMux
    port map (
            O => \N__39136\,
            I => \N__39131\
        );

    \I__7620\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39126\
        );

    \I__7619\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39126\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__39131\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_27\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__39126\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_27\
        );

    \I__7616\ : InMux
    port map (
            O => \N__39121\,
            I => \N__39115\
        );

    \I__7615\ : InMux
    port map (
            O => \N__39120\,
            I => \N__39115\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__39115\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\
        );

    \I__7613\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39107\
        );

    \I__7612\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39102\
        );

    \I__7611\ : InMux
    port map (
            O => \N__39110\,
            I => \N__39102\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__39107\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_26\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__39102\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_26\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__39097\,
            I => \N__39094\
        );

    \I__7607\ : InMux
    port map (
            O => \N__39094\,
            I => \N__39091\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__39091\,
            I => \N__39088\
        );

    \I__7605\ : Odrv12
    port map (
            O => \N__39088\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\
        );

    \I__7604\ : CascadeMux
    port map (
            O => \N__39085\,
            I => \N__39081\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__39084\,
            I => \N__39078\
        );

    \I__7602\ : InMux
    port map (
            O => \N__39081\,
            I => \N__39073\
        );

    \I__7601\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39073\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__39073\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\
        );

    \I__7599\ : InMux
    port map (
            O => \N__39070\,
            I => \bfn_14_11_0_\
        );

    \I__7598\ : InMux
    port map (
            O => \N__39067\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__7597\ : InMux
    port map (
            O => \N__39064\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__7596\ : InMux
    port map (
            O => \N__39061\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__7595\ : InMux
    port map (
            O => \N__39058\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__7594\ : InMux
    port map (
            O => \N__39055\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__7593\ : InMux
    port map (
            O => \N__39052\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__7592\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39044\
        );

    \I__7591\ : InMux
    port map (
            O => \N__39048\,
            I => \N__39039\
        );

    \I__7590\ : InMux
    port map (
            O => \N__39047\,
            I => \N__39039\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__39044\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_23\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__39039\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_23\
        );

    \I__7587\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39028\
        );

    \I__7586\ : InMux
    port map (
            O => \N__39033\,
            I => \N__39028\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__39028\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__39025\,
            I => \N__39020\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__39024\,
            I => \N__39017\
        );

    \I__7582\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39014\
        );

    \I__7581\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39009\
        );

    \I__7580\ : InMux
    port map (
            O => \N__39017\,
            I => \N__39009\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__39014\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_22\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__39009\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_22\
        );

    \I__7577\ : InMux
    port map (
            O => \N__39004\,
            I => \N__39001\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__39001\,
            I => \N__38998\
        );

    \I__7575\ : Odrv12
    port map (
            O => \N__38998\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\
        );

    \I__7574\ : InMux
    port map (
            O => \N__38995\,
            I => \N__38989\
        );

    \I__7573\ : InMux
    port map (
            O => \N__38994\,
            I => \N__38989\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__38989\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\
        );

    \I__7571\ : InMux
    port map (
            O => \N__38986\,
            I => \N__38983\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__38983\,
            I => \N__38980\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__38980\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt24\
        );

    \I__7568\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38971\
        );

    \I__7567\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38971\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__38971\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\
        );

    \I__7565\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38963\
        );

    \I__7564\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38958\
        );

    \I__7563\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38958\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__38963\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__38958\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_25\
        );

    \I__7560\ : CascadeMux
    port map (
            O => \N__38953\,
            I => \N__38948\
        );

    \I__7559\ : CascadeMux
    port map (
            O => \N__38952\,
            I => \N__38945\
        );

    \I__7558\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38942\
        );

    \I__7557\ : InMux
    port map (
            O => \N__38948\,
            I => \N__38937\
        );

    \I__7556\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38937\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__38942\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_24\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__38937\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_24\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__38932\,
            I => \N__38929\
        );

    \I__7552\ : InMux
    port map (
            O => \N__38929\,
            I => \N__38926\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38923\
        );

    \I__7550\ : Odrv4
    port map (
            O => \N__38923\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\
        );

    \I__7549\ : InMux
    port map (
            O => \N__38920\,
            I => \N__38914\
        );

    \I__7548\ : InMux
    port map (
            O => \N__38919\,
            I => \N__38914\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__38914\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\
        );

    \I__7546\ : InMux
    port map (
            O => \N__38911\,
            I => \N__38908\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__38908\,
            I => \N__38905\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__38905\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt26\
        );

    \I__7543\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38896\
        );

    \I__7542\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38896\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__38896\,
            I => \N__38893\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__38893\,
            I => \N__38890\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__38890\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__38887\,
            I => \N__38883\
        );

    \I__7537\ : InMux
    port map (
            O => \N__38886\,
            I => \N__38878\
        );

    \I__7536\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38878\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__38878\,
            I => \N__38875\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__38875\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__38872\,
            I => \N__38867\
        );

    \I__7532\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38864\
        );

    \I__7531\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38859\
        );

    \I__7530\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38859\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__38864\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_17\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__38859\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_17\
        );

    \I__7527\ : InMux
    port map (
            O => \N__38854\,
            I => \N__38849\
        );

    \I__7526\ : InMux
    port map (
            O => \N__38853\,
            I => \N__38844\
        );

    \I__7525\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38844\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__38849\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_16\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__38844\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_16\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__38839\,
            I => \N__38836\
        );

    \I__7521\ : InMux
    port map (
            O => \N__38836\,
            I => \N__38833\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__38833\,
            I => \N__38830\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__38830\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\
        );

    \I__7518\ : InMux
    port map (
            O => \N__38827\,
            I => \N__38824\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__38824\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__7516\ : CascadeMux
    port map (
            O => \N__38821\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\
        );

    \I__7515\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38813\
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__38817\,
            I => \N__38809\
        );

    \I__7513\ : InMux
    port map (
            O => \N__38816\,
            I => \N__38804\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__38813\,
            I => \N__38801\
        );

    \I__7511\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38798\
        );

    \I__7510\ : InMux
    port map (
            O => \N__38809\,
            I => \N__38791\
        );

    \I__7509\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38791\
        );

    \I__7508\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38791\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__38804\,
            I => \N__38786\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__38801\,
            I => \N__38786\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__38798\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__38791\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__38786\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7502\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38776\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__38776\,
            I => \N__38772\
        );

    \I__7500\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38769\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__38772\,
            I => \N__38764\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__38769\,
            I => \N__38764\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__38764\,
            I => \N__38760\
        );

    \I__7496\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38757\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__38760\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__38757\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__7493\ : CascadeMux
    port map (
            O => \N__38752\,
            I => \N__38748\
        );

    \I__7492\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38745\
        );

    \I__7491\ : InMux
    port map (
            O => \N__38748\,
            I => \N__38742\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__38745\,
            I => \phase_controller_inst1.stoper_hc.counter\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__38742\,
            I => \phase_controller_inst1.stoper_hc.counter\
        );

    \I__7488\ : InMux
    port map (
            O => \N__38737\,
            I => \N__38732\
        );

    \I__7487\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38727\
        );

    \I__7486\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38727\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__38732\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_21\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__38727\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_21\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__38722\,
            I => \N__38717\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__38721\,
            I => \N__38714\
        );

    \I__7481\ : InMux
    port map (
            O => \N__38720\,
            I => \N__38711\
        );

    \I__7480\ : InMux
    port map (
            O => \N__38717\,
            I => \N__38706\
        );

    \I__7479\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38706\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__38711\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_20\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__38706\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_20\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__38701\,
            I => \N__38698\
        );

    \I__7475\ : InMux
    port map (
            O => \N__38698\,
            I => \N__38695\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__38695\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt20\
        );

    \I__7473\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38686\
        );

    \I__7472\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38686\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__38686\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\
        );

    \I__7470\ : InMux
    port map (
            O => \N__38683\,
            I => \N__38677\
        );

    \I__7469\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38677\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__38677\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\
        );

    \I__7467\ : CascadeMux
    port map (
            O => \N__38674\,
            I => \N__38671\
        );

    \I__7466\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38668\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__38668\,
            I => \N__38665\
        );

    \I__7464\ : Odrv12
    port map (
            O => \N__38665\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt22\
        );

    \I__7463\ : InMux
    port map (
            O => \N__38662\,
            I => \N__38659\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__38659\,
            I => \N__38656\
        );

    \I__7461\ : Span4Mux_h
    port map (
            O => \N__38656\,
            I => \N__38653\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__38653\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt28\
        );

    \I__7459\ : CascadeMux
    port map (
            O => \N__38650\,
            I => \N__38647\
        );

    \I__7458\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38644\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__38644\,
            I => \N__38641\
        );

    \I__7456\ : Span12Mux_h
    port map (
            O => \N__38641\,
            I => \N__38638\
        );

    \I__7455\ : Odrv12
    port map (
            O => \N__38638\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\
        );

    \I__7454\ : InMux
    port map (
            O => \N__38635\,
            I => \N__38632\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__38632\,
            I => \N__38629\
        );

    \I__7452\ : Span4Mux_h
    port map (
            O => \N__38629\,
            I => \N__38626\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__38626\,
            I => \N__38623\
        );

    \I__7450\ : Odrv4
    port map (
            O => \N__38623\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt30\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__38620\,
            I => \N__38617\
        );

    \I__7448\ : InMux
    port map (
            O => \N__38617\,
            I => \N__38614\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__38614\,
            I => \N__38611\
        );

    \I__7446\ : Span4Mux_v
    port map (
            O => \N__38611\,
            I => \N__38608\
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__38608\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\
        );

    \I__7444\ : InMux
    port map (
            O => \N__38605\,
            I => \bfn_14_8_0_\
        );

    \I__7443\ : InMux
    port map (
            O => \N__38602\,
            I => \N__38599\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__38599\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\
        );

    \I__7441\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38593\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__38593\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt16\
        );

    \I__7439\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38587\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__38587\,
            I => \N__38583\
        );

    \I__7437\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38580\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__38583\,
            I => \N__38577\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__38580\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_10\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__38577\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_10\
        );

    \I__7433\ : CascadeMux
    port map (
            O => \N__38572\,
            I => \N__38569\
        );

    \I__7432\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38566\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__38566\,
            I => \phase_controller_inst1.stoper_hc.counter_i_10\
        );

    \I__7430\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38559\
        );

    \I__7429\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38556\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__38559\,
            I => \N__38553\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__38556\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_11\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__38553\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_11\
        );

    \I__7425\ : CascadeMux
    port map (
            O => \N__38548\,
            I => \N__38545\
        );

    \I__7424\ : InMux
    port map (
            O => \N__38545\,
            I => \N__38542\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__38542\,
            I => \phase_controller_inst1.stoper_hc.counter_i_11\
        );

    \I__7422\ : InMux
    port map (
            O => \N__38539\,
            I => \N__38535\
        );

    \I__7421\ : InMux
    port map (
            O => \N__38538\,
            I => \N__38532\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__38535\,
            I => \N__38529\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__38532\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_12\
        );

    \I__7418\ : Odrv4
    port map (
            O => \N__38529\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_12\
        );

    \I__7417\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38521\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__38521\,
            I => \phase_controller_inst1.stoper_hc.counter_i_12\
        );

    \I__7415\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38515\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__38515\,
            I => \N__38511\
        );

    \I__7413\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38508\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__38511\,
            I => \N__38505\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__38508\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_13\
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__38505\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_13\
        );

    \I__7409\ : CascadeMux
    port map (
            O => \N__38500\,
            I => \N__38497\
        );

    \I__7408\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38494\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__38494\,
            I => \N__38491\
        );

    \I__7406\ : Odrv4
    port map (
            O => \N__38491\,
            I => \phase_controller_inst1.stoper_hc.counter_i_13\
        );

    \I__7405\ : InMux
    port map (
            O => \N__38488\,
            I => \N__38484\
        );

    \I__7404\ : InMux
    port map (
            O => \N__38487\,
            I => \N__38481\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__38484\,
            I => \N__38478\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__38481\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_14\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__38478\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_14\
        );

    \I__7400\ : CascadeMux
    port map (
            O => \N__38473\,
            I => \N__38470\
        );

    \I__7399\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38467\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__38467\,
            I => \phase_controller_inst1.stoper_hc.counter_i_14\
        );

    \I__7397\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38461\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__38461\,
            I => \N__38457\
        );

    \I__7395\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38454\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__38457\,
            I => \N__38451\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__38454\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_15\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__38451\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_15\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__38446\,
            I => \N__38443\
        );

    \I__7390\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38440\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__38440\,
            I => \phase_controller_inst1.stoper_hc.counter_i_15\
        );

    \I__7388\ : InMux
    port map (
            O => \N__38437\,
            I => \N__38434\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__38434\,
            I => \phase_controller_inst1.stoper_hc.un6_running_lt18\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__38431\,
            I => \N__38428\
        );

    \I__7385\ : InMux
    port map (
            O => \N__38428\,
            I => \N__38425\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__38425\,
            I => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\
        );

    \I__7383\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38418\
        );

    \I__7382\ : InMux
    port map (
            O => \N__38421\,
            I => \N__38415\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__38418\,
            I => \N__38412\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__38415\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_2\
        );

    \I__7379\ : Odrv4
    port map (
            O => \N__38412\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_2\
        );

    \I__7378\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38404\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__38404\,
            I => \phase_controller_inst1.stoper_hc.counter_i_2\
        );

    \I__7376\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38398\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__38398\,
            I => \N__38394\
        );

    \I__7374\ : InMux
    port map (
            O => \N__38397\,
            I => \N__38391\
        );

    \I__7373\ : Span4Mux_v
    port map (
            O => \N__38394\,
            I => \N__38388\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__38391\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_3\
        );

    \I__7371\ : Odrv4
    port map (
            O => \N__38388\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_3\
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__38383\,
            I => \N__38380\
        );

    \I__7369\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38377\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__38377\,
            I => \phase_controller_inst1.stoper_hc.counter_i_3\
        );

    \I__7367\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38370\
        );

    \I__7366\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38367\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__38370\,
            I => \N__38364\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__38367\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_4\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__38364\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_4\
        );

    \I__7362\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38356\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__38356\,
            I => \phase_controller_inst1.stoper_hc.counter_i_4\
        );

    \I__7360\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38350\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__38350\,
            I => \N__38346\
        );

    \I__7358\ : InMux
    port map (
            O => \N__38349\,
            I => \N__38343\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__38346\,
            I => \N__38340\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__38343\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_5\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__38340\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_5\
        );

    \I__7354\ : CascadeMux
    port map (
            O => \N__38335\,
            I => \N__38332\
        );

    \I__7353\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38329\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__38329\,
            I => \phase_controller_inst1.stoper_hc.counter_i_5\
        );

    \I__7351\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38323\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__38323\,
            I => \N__38319\
        );

    \I__7349\ : InMux
    port map (
            O => \N__38322\,
            I => \N__38316\
        );

    \I__7348\ : Span4Mux_v
    port map (
            O => \N__38319\,
            I => \N__38313\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__38316\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_6\
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__38313\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_6\
        );

    \I__7345\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__38305\,
            I => \phase_controller_inst1.stoper_hc.counter_i_6\
        );

    \I__7343\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38298\
        );

    \I__7342\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38295\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38292\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__38295\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_7\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__38292\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_7\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__38287\,
            I => \N__38284\
        );

    \I__7337\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38281\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__38281\,
            I => \N__38278\
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__38278\,
            I => \phase_controller_inst1.stoper_hc.counter_i_7\
        );

    \I__7334\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__38272\,
            I => \N__38268\
        );

    \I__7332\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38265\
        );

    \I__7331\ : Span4Mux_h
    port map (
            O => \N__38268\,
            I => \N__38262\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__38265\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_8\
        );

    \I__7329\ : Odrv4
    port map (
            O => \N__38262\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_8\
        );

    \I__7328\ : CascadeMux
    port map (
            O => \N__38257\,
            I => \N__38254\
        );

    \I__7327\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38251\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__38251\,
            I => \phase_controller_inst1.stoper_hc.counter_i_8\
        );

    \I__7325\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38244\
        );

    \I__7324\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38241\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__38244\,
            I => \N__38238\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__38241\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_9\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__38238\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_9\
        );

    \I__7320\ : CascadeMux
    port map (
            O => \N__38233\,
            I => \N__38230\
        );

    \I__7319\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__38227\,
            I => \phase_controller_inst1.stoper_hc.counter_i_9\
        );

    \I__7317\ : InMux
    port map (
            O => \N__38224\,
            I => \N__38221\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__38221\,
            I => \N__38218\
        );

    \I__7315\ : Odrv4
    port map (
            O => \N__38218\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__7314\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38212\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__38212\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__7312\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38206\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__38206\,
            I => \N__38202\
        );

    \I__7310\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38199\
        );

    \I__7309\ : Span12Mux_v
    port map (
            O => \N__38202\,
            I => \N__38196\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__38199\,
            I => \N__38191\
        );

    \I__7307\ : Span12Mux_h
    port map (
            O => \N__38196\,
            I => \N__38191\
        );

    \I__7306\ : Odrv12
    port map (
            O => \N__38191\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__7305\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__38185\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__7303\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38178\
        );

    \I__7302\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38175\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__38178\,
            I => \N__38172\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__38175\,
            I => \N__38169\
        );

    \I__7299\ : Span12Mux_s10_v
    port map (
            O => \N__38172\,
            I => \N__38166\
        );

    \I__7298\ : Odrv4
    port map (
            O => \N__38169\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__7297\ : Odrv12
    port map (
            O => \N__38166\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__7296\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38158\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__38158\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__7294\ : CascadeMux
    port map (
            O => \N__38155\,
            I => \N__38151\
        );

    \I__7293\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38143\
        );

    \I__7292\ : InMux
    port map (
            O => \N__38151\,
            I => \N__38143\
        );

    \I__7291\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38143\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__38143\,
            I => \N__38140\
        );

    \I__7289\ : Odrv12
    port map (
            O => \N__38140\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7288\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38131\
        );

    \I__7287\ : InMux
    port map (
            O => \N__38136\,
            I => \N__38131\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__38131\,
            I => \N__38128\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__38128\,
            I => \N__38123\
        );

    \I__7284\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38118\
        );

    \I__7283\ : InMux
    port map (
            O => \N__38126\,
            I => \N__38118\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__38123\,
            I => \N__38115\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__38118\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__38115\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7279\ : ClkMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__7278\ : GlobalMux
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__7277\ : gio2CtrlBuf
    port map (
            O => \N__38104\,
            I => delay_tr_input_c_g
        );

    \I__7276\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38097\
        );

    \I__7275\ : CascadeMux
    port map (
            O => \N__38100\,
            I => \N__38092\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__38097\,
            I => \N__38089\
        );

    \I__7273\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38084\
        );

    \I__7272\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38084\
        );

    \I__7271\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38081\
        );

    \I__7270\ : Span12Mux_v
    port map (
            O => \N__38089\,
            I => \N__38078\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__38084\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__38081\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7267\ : Odrv12
    port map (
            O => \N__38078\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7266\ : IoInMux
    port map (
            O => \N__38071\,
            I => \N__38068\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__38068\,
            I => \N__38065\
        );

    \I__7264\ : Odrv12
    port map (
            O => \N__38065\,
            I => s2_phy_c
        );

    \I__7263\ : InMux
    port map (
            O => \N__38062\,
            I => \N__38059\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__38059\,
            I => \N__38055\
        );

    \I__7261\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38052\
        );

    \I__7260\ : Span4Mux_h
    port map (
            O => \N__38055\,
            I => \N__38049\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__38052\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_0\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__38049\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_0\
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__38044\,
            I => \N__38041\
        );

    \I__7256\ : InMux
    port map (
            O => \N__38041\,
            I => \N__38038\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__38038\,
            I => \phase_controller_inst1.stoper_hc.counter_i_0\
        );

    \I__7254\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38032\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__38032\,
            I => \N__38028\
        );

    \I__7252\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38025\
        );

    \I__7251\ : Span4Mux_h
    port map (
            O => \N__38028\,
            I => \N__38022\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__38025\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_1\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__38022\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_1\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__38017\,
            I => \N__38014\
        );

    \I__7247\ : InMux
    port map (
            O => \N__38014\,
            I => \N__38011\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__38011\,
            I => \phase_controller_inst1.stoper_hc.counter_i_1\
        );

    \I__7245\ : InMux
    port map (
            O => \N__38008\,
            I => \N__38005\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__38005\,
            I => \N__38001\
        );

    \I__7243\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37998\
        );

    \I__7242\ : Span4Mux_s2_h
    port map (
            O => \N__38001\,
            I => \N__37995\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__37998\,
            I => \N__37992\
        );

    \I__7240\ : Sp12to4
    port map (
            O => \N__37995\,
            I => \N__37989\
        );

    \I__7239\ : Span4Mux_v
    port map (
            O => \N__37992\,
            I => \N__37986\
        );

    \I__7238\ : Span12Mux_s11_v
    port map (
            O => \N__37989\,
            I => \N__37983\
        );

    \I__7237\ : Odrv4
    port map (
            O => \N__37986\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__7236\ : Odrv12
    port map (
            O => \N__37983\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__7235\ : CascadeMux
    port map (
            O => \N__37978\,
            I => \N__37975\
        );

    \I__7234\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37972\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__37972\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__7232\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37966\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__37963\,
            I => \N__37959\
        );

    \I__7229\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37956\
        );

    \I__7228\ : Sp12to4
    port map (
            O => \N__37959\,
            I => \N__37953\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__37956\,
            I => \N__37948\
        );

    \I__7226\ : Span12Mux_h
    port map (
            O => \N__37953\,
            I => \N__37948\
        );

    \I__7225\ : Odrv12
    port map (
            O => \N__37948\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__7224\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37942\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__37942\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__7222\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37935\
        );

    \I__7221\ : InMux
    port map (
            O => \N__37938\,
            I => \N__37932\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__37935\,
            I => \N__37929\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__37932\,
            I => \N__37926\
        );

    \I__7218\ : Span12Mux_s11_v
    port map (
            O => \N__37929\,
            I => \N__37923\
        );

    \I__7217\ : Odrv4
    port map (
            O => \N__37926\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__7216\ : Odrv12
    port map (
            O => \N__37923\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__7215\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37915\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__37915\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__7213\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37909\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__37909\,
            I => \N__37905\
        );

    \I__7211\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37902\
        );

    \I__7210\ : Span12Mux_s6_v
    port map (
            O => \N__37905\,
            I => \N__37899\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__37902\,
            I => \N__37896\
        );

    \I__7208\ : Span12Mux_h
    port map (
            O => \N__37899\,
            I => \N__37893\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__37896\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__7206\ : Odrv12
    port map (
            O => \N__37893\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__7205\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37885\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__37885\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__7203\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__37879\,
            I => \N__37875\
        );

    \I__7201\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37872\
        );

    \I__7200\ : Span12Mux_v
    port map (
            O => \N__37875\,
            I => \N__37869\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__37872\,
            I => \N__37864\
        );

    \I__7198\ : Span12Mux_h
    port map (
            O => \N__37869\,
            I => \N__37864\
        );

    \I__7197\ : Odrv12
    port map (
            O => \N__37864\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__7196\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37858\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__37858\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__7194\ : InMux
    port map (
            O => \N__37855\,
            I => \N__37852\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__37852\,
            I => \N__37849\
        );

    \I__7192\ : Span4Mux_s1_h
    port map (
            O => \N__37849\,
            I => \N__37845\
        );

    \I__7191\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37842\
        );

    \I__7190\ : Sp12to4
    port map (
            O => \N__37845\,
            I => \N__37839\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__37842\,
            I => \N__37836\
        );

    \I__7188\ : Span12Mux_s10_v
    port map (
            O => \N__37839\,
            I => \N__37833\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__37836\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__7186\ : Odrv12
    port map (
            O => \N__37833\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__7185\ : InMux
    port map (
            O => \N__37828\,
            I => \N__37825\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__37825\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__7183\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37818\
        );

    \I__7182\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37815\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__37818\,
            I => \N__37812\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__37815\,
            I => \N__37807\
        );

    \I__7179\ : Span12Mux_s7_v
    port map (
            O => \N__37812\,
            I => \N__37807\
        );

    \I__7178\ : Span12Mux_h
    port map (
            O => \N__37807\,
            I => \N__37804\
        );

    \I__7177\ : Odrv12
    port map (
            O => \N__37804\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__7176\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37798\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__37798\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__7174\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__37792\,
            I => \N__37789\
        );

    \I__7172\ : Sp12to4
    port map (
            O => \N__37789\,
            I => \N__37785\
        );

    \I__7171\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37782\
        );

    \I__7170\ : Span12Mux_v
    port map (
            O => \N__37785\,
            I => \N__37779\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__37782\,
            I => \N__37774\
        );

    \I__7168\ : Span12Mux_h
    port map (
            O => \N__37779\,
            I => \N__37774\
        );

    \I__7167\ : Odrv12
    port map (
            O => \N__37774\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__7166\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37768\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__37768\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__7164\ : InMux
    port map (
            O => \N__37765\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__7163\ : InMux
    port map (
            O => \N__37762\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__7162\ : InMux
    port map (
            O => \N__37759\,
            I => \N__37753\
        );

    \I__7161\ : InMux
    port map (
            O => \N__37758\,
            I => \N__37753\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__37753\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__7159\ : InMux
    port map (
            O => \N__37750\,
            I => \N__37744\
        );

    \I__7158\ : InMux
    port map (
            O => \N__37749\,
            I => \N__37744\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__37744\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__7156\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37735\
        );

    \I__7155\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37735\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__37735\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__37732\,
            I => \N__37728\
        );

    \I__7152\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37723\
        );

    \I__7151\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37723\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__37723\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__7149\ : CascadeMux
    port map (
            O => \N__37720\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__7148\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37714\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__37714\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__37711\,
            I => \N__37708\
        );

    \I__7145\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37705\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37700\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__37704\,
            I => \N__37697\
        );

    \I__7142\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37693\
        );

    \I__7141\ : Span4Mux_h
    port map (
            O => \N__37700\,
            I => \N__37690\
        );

    \I__7140\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37687\
        );

    \I__7139\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37684\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__37693\,
            I => \N__37681\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__37690\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__37687\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__37684\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__37681\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__7133\ : CascadeMux
    port map (
            O => \N__37672\,
            I => \N__37668\
        );

    \I__7132\ : InMux
    port map (
            O => \N__37671\,
            I => \N__37664\
        );

    \I__7131\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37661\
        );

    \I__7130\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37658\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37654\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__37661\,
            I => \N__37651\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__37658\,
            I => \N__37648\
        );

    \I__7126\ : InMux
    port map (
            O => \N__37657\,
            I => \N__37645\
        );

    \I__7125\ : Span4Mux_h
    port map (
            O => \N__37654\,
            I => \N__37642\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__37651\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7123\ : Odrv12
    port map (
            O => \N__37648\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__37645\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__37642\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__7120\ : CascadeMux
    port map (
            O => \N__37633\,
            I => \N__37629\
        );

    \I__7119\ : CascadeMux
    port map (
            O => \N__37632\,
            I => \N__37626\
        );

    \I__7118\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37623\
        );

    \I__7117\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37620\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__37623\,
            I => \N__37616\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37613\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__37619\,
            I => \N__37610\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__37616\,
            I => \N__37606\
        );

    \I__7112\ : Span4Mux_h
    port map (
            O => \N__37613\,
            I => \N__37603\
        );

    \I__7111\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37600\
        );

    \I__7110\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37597\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__37606\,
            I => \N__37594\
        );

    \I__7108\ : Odrv4
    port map (
            O => \N__37603\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__37600\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__37597\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7105\ : Odrv4
    port map (
            O => \N__37594\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__7104\ : InMux
    port map (
            O => \N__37585\,
            I => \N__37581\
        );

    \I__7103\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37576\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__37581\,
            I => \N__37573\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__37580\,
            I => \N__37570\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__37579\,
            I => \N__37567\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__37576\,
            I => \N__37564\
        );

    \I__7098\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37561\
        );

    \I__7097\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37558\
        );

    \I__7096\ : InMux
    port map (
            O => \N__37567\,
            I => \N__37555\
        );

    \I__7095\ : Span4Mux_h
    port map (
            O => \N__37564\,
            I => \N__37552\
        );

    \I__7094\ : Odrv4
    port map (
            O => \N__37561\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__37558\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__37555\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7091\ : Odrv4
    port map (
            O => \N__37552\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__7090\ : InMux
    port map (
            O => \N__37543\,
            I => \N__37540\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__37540\,
            I => \N__37537\
        );

    \I__7088\ : Span4Mux_h
    port map (
            O => \N__37537\,
            I => \N__37534\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__37534\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__7086\ : InMux
    port map (
            O => \N__37531\,
            I => \N__37528\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__37528\,
            I => \N__37524\
        );

    \I__7084\ : InMux
    port map (
            O => \N__37527\,
            I => \N__37521\
        );

    \I__7083\ : Span12Mux_v
    port map (
            O => \N__37524\,
            I => \N__37518\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__37521\,
            I => \N__37513\
        );

    \I__7081\ : Span12Mux_h
    port map (
            O => \N__37518\,
            I => \N__37513\
        );

    \I__7080\ : Odrv12
    port map (
            O => \N__37513\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__7079\ : InMux
    port map (
            O => \N__37510\,
            I => \N__37507\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__37507\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__7077\ : InMux
    port map (
            O => \N__37504\,
            I => \N__37501\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__37501\,
            I => \N__37498\
        );

    \I__7075\ : Span4Mux_s3_h
    port map (
            O => \N__37498\,
            I => \N__37494\
        );

    \I__7074\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37491\
        );

    \I__7073\ : Span4Mux_h
    port map (
            O => \N__37494\,
            I => \N__37488\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__37491\,
            I => \N__37483\
        );

    \I__7071\ : Span4Mux_h
    port map (
            O => \N__37488\,
            I => \N__37483\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__37483\,
            I => \N__37480\
        );

    \I__7069\ : Odrv4
    port map (
            O => \N__37480\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__7068\ : InMux
    port map (
            O => \N__37477\,
            I => \N__37474\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__37474\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__7066\ : InMux
    port map (
            O => \N__37471\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__7065\ : InMux
    port map (
            O => \N__37468\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__7064\ : InMux
    port map (
            O => \N__37465\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__7063\ : InMux
    port map (
            O => \N__37462\,
            I => \bfn_13_20_0_\
        );

    \I__7062\ : InMux
    port map (
            O => \N__37459\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__7061\ : InMux
    port map (
            O => \N__37456\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__7060\ : InMux
    port map (
            O => \N__37453\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__7059\ : InMux
    port map (
            O => \N__37450\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__7058\ : InMux
    port map (
            O => \N__37447\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__7057\ : InMux
    port map (
            O => \N__37444\,
            I => \N__37441\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__37441\,
            I => \N__37438\
        );

    \I__7055\ : Span4Mux_v
    port map (
            O => \N__37438\,
            I => \N__37435\
        );

    \I__7054\ : Sp12to4
    port map (
            O => \N__37435\,
            I => \N__37431\
        );

    \I__7053\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37428\
        );

    \I__7052\ : Span12Mux_h
    port map (
            O => \N__37431\,
            I => \N__37425\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__37428\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7050\ : Odrv12
    port map (
            O => \N__37425\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__7049\ : InMux
    port map (
            O => \N__37420\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__7048\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37414\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__37414\,
            I => \N__37411\
        );

    \I__7046\ : Span4Mux_v
    port map (
            O => \N__37411\,
            I => \N__37408\
        );

    \I__7045\ : Sp12to4
    port map (
            O => \N__37408\,
            I => \N__37405\
        );

    \I__7044\ : Span12Mux_h
    port map (
            O => \N__37405\,
            I => \N__37401\
        );

    \I__7043\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37398\
        );

    \I__7042\ : Span12Mux_v
    port map (
            O => \N__37401\,
            I => \N__37395\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__37398\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7040\ : Odrv12
    port map (
            O => \N__37395\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__7039\ : InMux
    port map (
            O => \N__37390\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37384\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__37384\,
            I => \N__37381\
        );

    \I__7036\ : Span4Mux_v
    port map (
            O => \N__37381\,
            I => \N__37378\
        );

    \I__7035\ : Sp12to4
    port map (
            O => \N__37378\,
            I => \N__37375\
        );

    \I__7034\ : Span12Mux_s11_h
    port map (
            O => \N__37375\,
            I => \N__37371\
        );

    \I__7033\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37368\
        );

    \I__7032\ : Span12Mux_v
    port map (
            O => \N__37371\,
            I => \N__37365\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__37368\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7030\ : Odrv12
    port map (
            O => \N__37365\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__7029\ : InMux
    port map (
            O => \N__37360\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__7028\ : InMux
    port map (
            O => \N__37357\,
            I => \N__37354\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__37354\,
            I => \N__37351\
        );

    \I__7026\ : Sp12to4
    port map (
            O => \N__37351\,
            I => \N__37347\
        );

    \I__7025\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37344\
        );

    \I__7024\ : Span12Mux_h
    port map (
            O => \N__37347\,
            I => \N__37341\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__37344\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__7022\ : Odrv12
    port map (
            O => \N__37341\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__7021\ : InMux
    port map (
            O => \N__37336\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__7020\ : InMux
    port map (
            O => \N__37333\,
            I => \N__37330\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__37330\,
            I => \N__37327\
        );

    \I__7018\ : Sp12to4
    port map (
            O => \N__37327\,
            I => \N__37324\
        );

    \I__7017\ : Span12Mux_v
    port map (
            O => \N__37324\,
            I => \N__37320\
        );

    \I__7016\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37317\
        );

    \I__7015\ : Span12Mux_h
    port map (
            O => \N__37320\,
            I => \N__37314\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__37317\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7013\ : Odrv12
    port map (
            O => \N__37314\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__7012\ : InMux
    port map (
            O => \N__37309\,
            I => \bfn_13_19_0_\
        );

    \I__7011\ : InMux
    port map (
            O => \N__37306\,
            I => \N__37303\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__37303\,
            I => \N__37300\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__37300\,
            I => \N__37297\
        );

    \I__7008\ : Sp12to4
    port map (
            O => \N__37297\,
            I => \N__37293\
        );

    \I__7007\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37290\
        );

    \I__7006\ : Span12Mux_h
    port map (
            O => \N__37293\,
            I => \N__37287\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__37290\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__7004\ : Odrv12
    port map (
            O => \N__37287\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__7003\ : InMux
    port map (
            O => \N__37282\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__7002\ : InMux
    port map (
            O => \N__37279\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__7001\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37273\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__37273\,
            I => \N__37270\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__37270\,
            I => \N__37267\
        );

    \I__6998\ : Span4Mux_h
    port map (
            O => \N__37267\,
            I => \N__37264\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__37264\,
            I => \N__37260\
        );

    \I__6996\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37257\
        );

    \I__6995\ : Span4Mux_h
    port map (
            O => \N__37260\,
            I => \N__37254\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__37257\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__37254\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__6992\ : InMux
    port map (
            O => \N__37249\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__6991\ : InMux
    port map (
            O => \N__37246\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__6990\ : InMux
    port map (
            O => \N__37243\,
            I => \N__37240\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__37240\,
            I => \N__37237\
        );

    \I__6988\ : Sp12to4
    port map (
            O => \N__37237\,
            I => \N__37234\
        );

    \I__6987\ : Span12Mux_v
    port map (
            O => \N__37234\,
            I => \N__37230\
        );

    \I__6986\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37227\
        );

    \I__6985\ : Span12Mux_h
    port map (
            O => \N__37230\,
            I => \N__37224\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__37227\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__6983\ : Odrv12
    port map (
            O => \N__37224\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__6982\ : InMux
    port map (
            O => \N__37219\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__6981\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37213\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__37213\,
            I => \N__37210\
        );

    \I__6979\ : Sp12to4
    port map (
            O => \N__37210\,
            I => \N__37207\
        );

    \I__6978\ : Span12Mux_s9_v
    port map (
            O => \N__37207\,
            I => \N__37203\
        );

    \I__6977\ : InMux
    port map (
            O => \N__37206\,
            I => \N__37200\
        );

    \I__6976\ : Span12Mux_h
    port map (
            O => \N__37203\,
            I => \N__37197\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__37200\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__6974\ : Odrv12
    port map (
            O => \N__37197\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__6973\ : InMux
    port map (
            O => \N__37192\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__6972\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37186\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__37186\,
            I => \N__37183\
        );

    \I__6970\ : Sp12to4
    port map (
            O => \N__37183\,
            I => \N__37180\
        );

    \I__6969\ : Span12Mux_s10_v
    port map (
            O => \N__37180\,
            I => \N__37176\
        );

    \I__6968\ : InMux
    port map (
            O => \N__37179\,
            I => \N__37173\
        );

    \I__6967\ : Span12Mux_h
    port map (
            O => \N__37176\,
            I => \N__37170\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__37173\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6965\ : Odrv12
    port map (
            O => \N__37170\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6964\ : InMux
    port map (
            O => \N__37165\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__6963\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37159\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__37159\,
            I => \N__37156\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__37156\,
            I => \N__37153\
        );

    \I__6960\ : Sp12to4
    port map (
            O => \N__37153\,
            I => \N__37149\
        );

    \I__6959\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37146\
        );

    \I__6958\ : Span12Mux_s10_h
    port map (
            O => \N__37149\,
            I => \N__37143\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__37146\,
            I => \N__37140\
        );

    \I__6956\ : Span12Mux_v
    port map (
            O => \N__37143\,
            I => \N__37137\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__37140\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6954\ : Odrv12
    port map (
            O => \N__37137\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__6953\ : InMux
    port map (
            O => \N__37132\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__6952\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37126\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__37126\,
            I => \N__37123\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__37123\,
            I => \N__37120\
        );

    \I__6949\ : Sp12to4
    port map (
            O => \N__37120\,
            I => \N__37116\
        );

    \I__6948\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37113\
        );

    \I__6947\ : Span12Mux_h
    port map (
            O => \N__37116\,
            I => \N__37110\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__37113\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6945\ : Odrv12
    port map (
            O => \N__37110\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6944\ : InMux
    port map (
            O => \N__37105\,
            I => \bfn_13_18_0_\
        );

    \I__6943\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37099\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__37099\,
            I => \N__37096\
        );

    \I__6941\ : Span12Mux_s1_h
    port map (
            O => \N__37096\,
            I => \N__37092\
        );

    \I__6940\ : InMux
    port map (
            O => \N__37095\,
            I => \N__37089\
        );

    \I__6939\ : Span12Mux_h
    port map (
            O => \N__37092\,
            I => \N__37086\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__37089\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6937\ : Odrv12
    port map (
            O => \N__37086\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__6936\ : InMux
    port map (
            O => \N__37081\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__6935\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37075\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__37075\,
            I => \N__37072\
        );

    \I__6933\ : Sp12to4
    port map (
            O => \N__37072\,
            I => \N__37069\
        );

    \I__6932\ : Span12Mux_s7_v
    port map (
            O => \N__37069\,
            I => \N__37065\
        );

    \I__6931\ : InMux
    port map (
            O => \N__37068\,
            I => \N__37062\
        );

    \I__6930\ : Span12Mux_h
    port map (
            O => \N__37065\,
            I => \N__37059\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__37062\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6928\ : Odrv12
    port map (
            O => \N__37059\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__6927\ : InMux
    port map (
            O => \N__37054\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__6926\ : InMux
    port map (
            O => \N__37051\,
            I => \N__37048\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__37048\,
            I => \N__37045\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__37045\,
            I => \N__37042\
        );

    \I__6923\ : Sp12to4
    port map (
            O => \N__37042\,
            I => \N__37038\
        );

    \I__6922\ : InMux
    port map (
            O => \N__37041\,
            I => \N__37035\
        );

    \I__6921\ : Span12Mux_h
    port map (
            O => \N__37038\,
            I => \N__37032\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__37035\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__6919\ : Odrv12
    port map (
            O => \N__37032\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__6918\ : InMux
    port map (
            O => \N__37027\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__6917\ : InMux
    port map (
            O => \N__37024\,
            I => \N__37021\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__37021\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__6915\ : InMux
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__37015\,
            I => \N__37012\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__37012\,
            I => \N__37009\
        );

    \I__6912\ : Sp12to4
    port map (
            O => \N__37009\,
            I => \N__37005\
        );

    \I__6911\ : InMux
    port map (
            O => \N__37008\,
            I => \N__37002\
        );

    \I__6910\ : Span12Mux_h
    port map (
            O => \N__37005\,
            I => \N__36999\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__37002\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6908\ : Odrv12
    port map (
            O => \N__36999\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__6907\ : InMux
    port map (
            O => \N__36994\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__6906\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36988\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__36988\,
            I => \N__36985\
        );

    \I__6904\ : Span12Mux_s1_h
    port map (
            O => \N__36985\,
            I => \N__36981\
        );

    \I__6903\ : InMux
    port map (
            O => \N__36984\,
            I => \N__36978\
        );

    \I__6902\ : Span12Mux_h
    port map (
            O => \N__36981\,
            I => \N__36975\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__36978\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6900\ : Odrv12
    port map (
            O => \N__36975\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__6899\ : InMux
    port map (
            O => \N__36970\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__6898\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36964\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__36964\,
            I => \N__36961\
        );

    \I__6896\ : Sp12to4
    port map (
            O => \N__36961\,
            I => \N__36958\
        );

    \I__6895\ : Span12Mux_s7_v
    port map (
            O => \N__36958\,
            I => \N__36954\
        );

    \I__6894\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36951\
        );

    \I__6893\ : Span12Mux_h
    port map (
            O => \N__36954\,
            I => \N__36948\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__36951\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6891\ : Odrv12
    port map (
            O => \N__36948\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__6890\ : InMux
    port map (
            O => \N__36943\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__6889\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36900\
        );

    \I__6888\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36900\
        );

    \I__6887\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36900\
        );

    \I__6886\ : InMux
    port map (
            O => \N__36937\,
            I => \N__36900\
        );

    \I__6885\ : InMux
    port map (
            O => \N__36936\,
            I => \N__36891\
        );

    \I__6884\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36891\
        );

    \I__6883\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36891\
        );

    \I__6882\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36891\
        );

    \I__6881\ : InMux
    port map (
            O => \N__36932\,
            I => \N__36882\
        );

    \I__6880\ : InMux
    port map (
            O => \N__36931\,
            I => \N__36882\
        );

    \I__6879\ : InMux
    port map (
            O => \N__36930\,
            I => \N__36882\
        );

    \I__6878\ : InMux
    port map (
            O => \N__36929\,
            I => \N__36882\
        );

    \I__6877\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36875\
        );

    \I__6876\ : InMux
    port map (
            O => \N__36927\,
            I => \N__36875\
        );

    \I__6875\ : InMux
    port map (
            O => \N__36926\,
            I => \N__36875\
        );

    \I__6874\ : InMux
    port map (
            O => \N__36925\,
            I => \N__36866\
        );

    \I__6873\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36866\
        );

    \I__6872\ : InMux
    port map (
            O => \N__36923\,
            I => \N__36866\
        );

    \I__6871\ : InMux
    port map (
            O => \N__36922\,
            I => \N__36866\
        );

    \I__6870\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36857\
        );

    \I__6869\ : InMux
    port map (
            O => \N__36920\,
            I => \N__36857\
        );

    \I__6868\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36857\
        );

    \I__6867\ : InMux
    port map (
            O => \N__36918\,
            I => \N__36857\
        );

    \I__6866\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36848\
        );

    \I__6865\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36848\
        );

    \I__6864\ : InMux
    port map (
            O => \N__36915\,
            I => \N__36848\
        );

    \I__6863\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36848\
        );

    \I__6862\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36837\
        );

    \I__6861\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36837\
        );

    \I__6860\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36837\
        );

    \I__6859\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36837\
        );

    \I__6858\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36837\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__36900\,
            I => \N__36820\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__36891\,
            I => \N__36820\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__36882\,
            I => \N__36820\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__36875\,
            I => \N__36820\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__36866\,
            I => \N__36820\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__36857\,
            I => \N__36820\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__36848\,
            I => \N__36820\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__36837\,
            I => \N__36820\
        );

    \I__6849\ : Odrv12
    port map (
            O => \N__36820\,
            I => \phase_controller_inst1.stoper_hc.start_latched_i_0\
        );

    \I__6848\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36807\
        );

    \I__6847\ : InMux
    port map (
            O => \N__36816\,
            I => \N__36807\
        );

    \I__6846\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36807\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__36814\,
            I => \N__36804\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__36807\,
            I => \N__36799\
        );

    \I__6843\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36794\
        );

    \I__6842\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36794\
        );

    \I__6841\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36791\
        );

    \I__6840\ : Span4Mux_h
    port map (
            O => \N__36799\,
            I => \N__36788\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__36794\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__36791\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__36788\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6836\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36777\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__36780\,
            I => \N__36773\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__36777\,
            I => \N__36767\
        );

    \I__6833\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36764\
        );

    \I__6832\ : InMux
    port map (
            O => \N__36773\,
            I => \N__36757\
        );

    \I__6831\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36757\
        );

    \I__6830\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36757\
        );

    \I__6829\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36754\
        );

    \I__6828\ : Span4Mux_h
    port map (
            O => \N__36767\,
            I => \N__36751\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__36764\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__36757\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__36754\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__36751\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__36742\,
            I => \N__36737\
        );

    \I__6822\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36734\
        );

    \I__6821\ : InMux
    port map (
            O => \N__36740\,
            I => \N__36731\
        );

    \I__6820\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36728\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__36734\,
            I => \N__36725\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__36731\,
            I => \N__36720\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__36728\,
            I => \N__36720\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__36725\,
            I => \N__36717\
        );

    \I__6815\ : Span4Mux_v
    port map (
            O => \N__36720\,
            I => \N__36714\
        );

    \I__6814\ : Span4Mux_h
    port map (
            O => \N__36717\,
            I => \N__36711\
        );

    \I__6813\ : Sp12to4
    port map (
            O => \N__36714\,
            I => \N__36708\
        );

    \I__6812\ : Odrv4
    port map (
            O => \N__36711\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\
        );

    \I__6811\ : Odrv12
    port map (
            O => \N__36708\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\
        );

    \I__6810\ : InMux
    port map (
            O => \N__36703\,
            I => \N__36700\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__36700\,
            I => \N__36696\
        );

    \I__6808\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36693\
        );

    \I__6807\ : Span4Mux_v
    port map (
            O => \N__36696\,
            I => \N__36687\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36684\
        );

    \I__6805\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36681\
        );

    \I__6804\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36678\
        );

    \I__6803\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36674\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__36687\,
            I => \N__36669\
        );

    \I__6801\ : Span4Mux_h
    port map (
            O => \N__36684\,
            I => \N__36669\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36666\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36663\
        );

    \I__6798\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36660\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__36674\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__36669\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__36666\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6794\ : Odrv4
    port map (
            O => \N__36663\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__36660\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__6792\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36646\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__36646\,
            I => \N__36643\
        );

    \I__6790\ : Span4Mux_h
    port map (
            O => \N__36643\,
            I => \N__36640\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__36640\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\
        );

    \I__6788\ : CEMux
    port map (
            O => \N__36637\,
            I => \N__36633\
        );

    \I__6787\ : CEMux
    port map (
            O => \N__36636\,
            I => \N__36630\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__36633\,
            I => \N__36625\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__36630\,
            I => \N__36625\
        );

    \I__6784\ : Span4Mux_v
    port map (
            O => \N__36625\,
            I => \N__36621\
        );

    \I__6783\ : CEMux
    port map (
            O => \N__36624\,
            I => \N__36618\
        );

    \I__6782\ : Span4Mux_h
    port map (
            O => \N__36621\,
            I => \N__36611\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__36618\,
            I => \N__36611\
        );

    \I__6780\ : CEMux
    port map (
            O => \N__36617\,
            I => \N__36608\
        );

    \I__6779\ : CEMux
    port map (
            O => \N__36616\,
            I => \N__36605\
        );

    \I__6778\ : Span4Mux_h
    port map (
            O => \N__36611\,
            I => \N__36602\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__36608\,
            I => \N__36599\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36596\
        );

    \I__6775\ : Sp12to4
    port map (
            O => \N__36602\,
            I => \N__36588\
        );

    \I__6774\ : Span12Mux_h
    port map (
            O => \N__36599\,
            I => \N__36588\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__36596\,
            I => \N__36585\
        );

    \I__6772\ : CEMux
    port map (
            O => \N__36595\,
            I => \N__36582\
        );

    \I__6771\ : CEMux
    port map (
            O => \N__36594\,
            I => \N__36579\
        );

    \I__6770\ : CEMux
    port map (
            O => \N__36593\,
            I => \N__36576\
        );

    \I__6769\ : Odrv12
    port map (
            O => \N__36588\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__36585\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__36582\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__36579\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__36576\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__6764\ : CEMux
    port map (
            O => \N__36565\,
            I => \N__36561\
        );

    \I__6763\ : CEMux
    port map (
            O => \N__36564\,
            I => \N__36558\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__36561\,
            I => \N__36553\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__36558\,
            I => \N__36550\
        );

    \I__6760\ : CEMux
    port map (
            O => \N__36557\,
            I => \N__36547\
        );

    \I__6759\ : CEMux
    port map (
            O => \N__36556\,
            I => \N__36544\
        );

    \I__6758\ : Span4Mux_v
    port map (
            O => \N__36553\,
            I => \N__36541\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__36550\,
            I => \N__36538\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__36547\,
            I => \N__36535\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__36544\,
            I => \N__36532\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__36541\,
            I => \N__36529\
        );

    \I__6753\ : Span4Mux_v
    port map (
            O => \N__36538\,
            I => \N__36526\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__36535\,
            I => \N__36523\
        );

    \I__6751\ : Span4Mux_h
    port map (
            O => \N__36532\,
            I => \N__36520\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__36529\,
            I => \N__36515\
        );

    \I__6749\ : Span4Mux_h
    port map (
            O => \N__36526\,
            I => \N__36515\
        );

    \I__6748\ : Span4Mux_h
    port map (
            O => \N__36523\,
            I => \N__36512\
        );

    \I__6747\ : Span4Mux_h
    port map (
            O => \N__36520\,
            I => \N__36509\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__36515\,
            I => \delay_measurement_inst.delay_tr_timer.N_168_i\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__36512\,
            I => \delay_measurement_inst.delay_tr_timer.N_168_i\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__36509\,
            I => \delay_measurement_inst.delay_tr_timer.N_168_i\
        );

    \I__6743\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36499\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__36499\,
            I => \N__36493\
        );

    \I__6741\ : InMux
    port map (
            O => \N__36498\,
            I => \N__36486\
        );

    \I__6740\ : InMux
    port map (
            O => \N__36497\,
            I => \N__36486\
        );

    \I__6739\ : InMux
    port map (
            O => \N__36496\,
            I => \N__36486\
        );

    \I__6738\ : Span4Mux_h
    port map (
            O => \N__36493\,
            I => \N__36483\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__36486\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__36483\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__6735\ : CEMux
    port map (
            O => \N__36478\,
            I => \N__36472\
        );

    \I__6734\ : CEMux
    port map (
            O => \N__36477\,
            I => \N__36469\
        );

    \I__6733\ : CEMux
    port map (
            O => \N__36476\,
            I => \N__36466\
        );

    \I__6732\ : CEMux
    port map (
            O => \N__36475\,
            I => \N__36463\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__36472\,
            I => \N__36459\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__36469\,
            I => \N__36456\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__36466\,
            I => \N__36453\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__36463\,
            I => \N__36450\
        );

    \I__6727\ : CEMux
    port map (
            O => \N__36462\,
            I => \N__36447\
        );

    \I__6726\ : Span4Mux_v
    port map (
            O => \N__36459\,
            I => \N__36444\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__36456\,
            I => \N__36441\
        );

    \I__6724\ : Span4Mux_v
    port map (
            O => \N__36453\,
            I => \N__36438\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__36450\,
            I => \N__36435\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36432\
        );

    \I__6721\ : Span4Mux_h
    port map (
            O => \N__36444\,
            I => \N__36429\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__36441\,
            I => \N__36426\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__36438\,
            I => \N__36421\
        );

    \I__6718\ : Span4Mux_h
    port map (
            O => \N__36435\,
            I => \N__36421\
        );

    \I__6717\ : Span4Mux_h
    port map (
            O => \N__36432\,
            I => \N__36418\
        );

    \I__6716\ : Odrv4
    port map (
            O => \N__36429\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__36426\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__36421\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__6713\ : Odrv4
    port map (
            O => \N__36418\,
            I => \delay_measurement_inst.delay_tr_timer.N_167_i\
        );

    \I__6712\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36406\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__36406\,
            I => \N__36401\
        );

    \I__6710\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36398\
        );

    \I__6709\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36395\
        );

    \I__6708\ : Span4Mux_v
    port map (
            O => \N__36401\,
            I => \N__36388\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__36398\,
            I => \N__36388\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__36395\,
            I => \N__36388\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__36388\,
            I => \N__36385\
        );

    \I__6704\ : Sp12to4
    port map (
            O => \N__36385\,
            I => \N__36382\
        );

    \I__6703\ : Span12Mux_h
    port map (
            O => \N__36382\,
            I => \N__36379\
        );

    \I__6702\ : Odrv12
    port map (
            O => \N__36379\,
            I => il_max_comp1_c
        );

    \I__6701\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36371\
        );

    \I__6700\ : InMux
    port map (
            O => \N__36375\,
            I => \N__36366\
        );

    \I__6699\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36366\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__36371\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__36366\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__6696\ : CascadeMux
    port map (
            O => \N__36361\,
            I => \phase_controller_inst1.stoper_hc.un4_start_0_cascade_\
        );

    \I__6695\ : InMux
    port map (
            O => \N__36358\,
            I => \N__36346\
        );

    \I__6694\ : InMux
    port map (
            O => \N__36357\,
            I => \N__36346\
        );

    \I__6693\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36346\
        );

    \I__6692\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36339\
        );

    \I__6691\ : InMux
    port map (
            O => \N__36354\,
            I => \N__36339\
        );

    \I__6690\ : InMux
    port map (
            O => \N__36353\,
            I => \N__36339\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__36346\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__36339\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__6687\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36329\
        );

    \I__6686\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36324\
        );

    \I__6685\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36324\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__36329\,
            I => \N__36321\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__36324\,
            I => \N__36318\
        );

    \I__6682\ : Span4Mux_v
    port map (
            O => \N__36321\,
            I => \N__36315\
        );

    \I__6681\ : Span4Mux_v
    port map (
            O => \N__36318\,
            I => \N__36312\
        );

    \I__6680\ : Sp12to4
    port map (
            O => \N__36315\,
            I => \N__36307\
        );

    \I__6679\ : Sp12to4
    port map (
            O => \N__36312\,
            I => \N__36307\
        );

    \I__6678\ : Span12Mux_h
    port map (
            O => \N__36307\,
            I => \N__36304\
        );

    \I__6677\ : Odrv12
    port map (
            O => \N__36304\,
            I => il_min_comp1_c
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__36301\,
            I => \N__36297\
        );

    \I__6675\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36294\
        );

    \I__6674\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36289\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36286\
        );

    \I__6672\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36281\
        );

    \I__6671\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36281\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__36289\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__36286\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__36281\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6667\ : CascadeMux
    port map (
            O => \N__36274\,
            I => \N__36269\
        );

    \I__6666\ : InMux
    port map (
            O => \N__36273\,
            I => \N__36265\
        );

    \I__6665\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36262\
        );

    \I__6664\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36257\
        );

    \I__6663\ : InMux
    port map (
            O => \N__36268\,
            I => \N__36257\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__36265\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__36262\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__36257\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6659\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__6658\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36244\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__36244\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__6656\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36238\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__36238\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__36235\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__6653\ : InMux
    port map (
            O => \N__36232\,
            I => \N__36229\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__36229\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__36226\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\
        );

    \I__6650\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36220\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__36220\,
            I => \N__36217\
        );

    \I__6648\ : Odrv4
    port map (
            O => \N__36217\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__6647\ : CEMux
    port map (
            O => \N__36214\,
            I => \N__36210\
        );

    \I__6646\ : CEMux
    port map (
            O => \N__36213\,
            I => \N__36206\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__36210\,
            I => \N__36202\
        );

    \I__6644\ : CEMux
    port map (
            O => \N__36209\,
            I => \N__36199\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__36206\,
            I => \N__36196\
        );

    \I__6642\ : CEMux
    port map (
            O => \N__36205\,
            I => \N__36193\
        );

    \I__6641\ : Span4Mux_v
    port map (
            O => \N__36202\,
            I => \N__36190\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__36187\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__36196\,
            I => \N__36184\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__36193\,
            I => \N__36181\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__36190\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6636\ : Odrv12
    port map (
            O => \N__36187\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6635\ : Odrv4
    port map (
            O => \N__36184\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6634\ : Odrv4
    port map (
            O => \N__36181\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6633\ : InMux
    port map (
            O => \N__36172\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_25\
        );

    \I__6632\ : InMux
    port map (
            O => \N__36169\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_26\
        );

    \I__6631\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36161\
        );

    \I__6630\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36156\
        );

    \I__6629\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36156\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__36161\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_28\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__36156\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_28\
        );

    \I__6626\ : InMux
    port map (
            O => \N__36151\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_27\
        );

    \I__6625\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36143\
        );

    \I__6624\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36138\
        );

    \I__6623\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36138\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__36143\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_29\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__36138\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_29\
        );

    \I__6620\ : InMux
    port map (
            O => \N__36133\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_28\
        );

    \I__6619\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36125\
        );

    \I__6618\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36122\
        );

    \I__6617\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36119\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__36125\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__36122\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__36119\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_30\
        );

    \I__6613\ : InMux
    port map (
            O => \N__36112\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_29\
        );

    \I__6612\ : InMux
    port map (
            O => \N__36109\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_30\
        );

    \I__6611\ : InMux
    port map (
            O => \N__36106\,
            I => \N__36101\
        );

    \I__6610\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36096\
        );

    \I__6609\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36096\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__36101\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__36096\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_31\
        );

    \I__6606\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36088\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__36088\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__6604\ : CascadeMux
    port map (
            O => \N__36085\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25_cascade_\
        );

    \I__6603\ : InMux
    port map (
            O => \N__36082\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_16\
        );

    \I__6602\ : InMux
    port map (
            O => \N__36079\,
            I => \N__36072\
        );

    \I__6601\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36072\
        );

    \I__6600\ : InMux
    port map (
            O => \N__36077\,
            I => \N__36069\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__36072\,
            I => \N__36066\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__36069\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_18\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__36066\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_18\
        );

    \I__6596\ : InMux
    port map (
            O => \N__36061\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_17\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__36058\,
            I => \N__36054\
        );

    \I__6594\ : CascadeMux
    port map (
            O => \N__36057\,
            I => \N__36051\
        );

    \I__6593\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36046\
        );

    \I__6592\ : InMux
    port map (
            O => \N__36051\,
            I => \N__36046\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36042\
        );

    \I__6590\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36039\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__36042\,
            I => \N__36036\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__36039\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_19\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__36036\,
            I => \phase_controller_inst1.stoper_hc.counterZ0Z_19\
        );

    \I__6586\ : InMux
    port map (
            O => \N__36031\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_18\
        );

    \I__6585\ : InMux
    port map (
            O => \N__36028\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_19\
        );

    \I__6584\ : InMux
    port map (
            O => \N__36025\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_20\
        );

    \I__6583\ : InMux
    port map (
            O => \N__36022\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_21\
        );

    \I__6582\ : InMux
    port map (
            O => \N__36019\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_22\
        );

    \I__6581\ : InMux
    port map (
            O => \N__36016\,
            I => \bfn_13_10_0_\
        );

    \I__6580\ : InMux
    port map (
            O => \N__36013\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_24\
        );

    \I__6579\ : InMux
    port map (
            O => \N__36010\,
            I => \bfn_13_8_0_\
        );

    \I__6578\ : InMux
    port map (
            O => \N__36007\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_8\
        );

    \I__6577\ : InMux
    port map (
            O => \N__36004\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_9\
        );

    \I__6576\ : InMux
    port map (
            O => \N__36001\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_10\
        );

    \I__6575\ : InMux
    port map (
            O => \N__35998\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_11\
        );

    \I__6574\ : InMux
    port map (
            O => \N__35995\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_12\
        );

    \I__6573\ : InMux
    port map (
            O => \N__35992\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_13\
        );

    \I__6572\ : InMux
    port map (
            O => \N__35989\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_14\
        );

    \I__6571\ : InMux
    port map (
            O => \N__35986\,
            I => \bfn_13_9_0_\
        );

    \I__6570\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35977\
        );

    \I__6569\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35977\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__35977\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\
        );

    \I__6567\ : InMux
    port map (
            O => \N__35974\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_0\
        );

    \I__6566\ : InMux
    port map (
            O => \N__35971\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_1\
        );

    \I__6565\ : InMux
    port map (
            O => \N__35968\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_2\
        );

    \I__6564\ : InMux
    port map (
            O => \N__35965\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_3\
        );

    \I__6563\ : InMux
    port map (
            O => \N__35962\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_4\
        );

    \I__6562\ : InMux
    port map (
            O => \N__35959\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_5\
        );

    \I__6561\ : InMux
    port map (
            O => \N__35956\,
            I => \phase_controller_inst1.stoper_hc.counter_cry_6\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__35953\,
            I => \N__35949\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__35952\,
            I => \N__35946\
        );

    \I__6558\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35943\
        );

    \I__6557\ : InMux
    port map (
            O => \N__35946\,
            I => \N__35939\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__35943\,
            I => \N__35936\
        );

    \I__6555\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35933\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__35939\,
            I => \N__35929\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__35936\,
            I => \N__35926\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__35933\,
            I => \N__35923\
        );

    \I__6551\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35920\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__35929\,
            I => \N__35913\
        );

    \I__6549\ : Span4Mux_h
    port map (
            O => \N__35926\,
            I => \N__35913\
        );

    \I__6548\ : Span4Mux_v
    port map (
            O => \N__35923\,
            I => \N__35913\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__35920\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__35913\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__6545\ : InMux
    port map (
            O => \N__35908\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__35905\,
            I => \N__35902\
        );

    \I__6543\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35899\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__35899\,
            I => \N__35894\
        );

    \I__6541\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35890\
        );

    \I__6540\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35887\
        );

    \I__6539\ : Span4Mux_v
    port map (
            O => \N__35894\,
            I => \N__35884\
        );

    \I__6538\ : InMux
    port map (
            O => \N__35893\,
            I => \N__35881\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__35890\,
            I => \N__35876\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__35887\,
            I => \N__35876\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__35884\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__35881\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__35876\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__6532\ : InMux
    port map (
            O => \N__35869\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__6531\ : InMux
    port map (
            O => \N__35866\,
            I => \N__35852\
        );

    \I__6530\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35845\
        );

    \I__6529\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35845\
        );

    \I__6528\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35845\
        );

    \I__6527\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35842\
        );

    \I__6526\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35833\
        );

    \I__6525\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35833\
        );

    \I__6524\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35833\
        );

    \I__6523\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35833\
        );

    \I__6522\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35830\
        );

    \I__6521\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35806\
        );

    \I__6520\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35806\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__35852\,
            I => \N__35803\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__35845\,
            I => \N__35800\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__35842\,
            I => \N__35797\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__35833\,
            I => \N__35792\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__35830\,
            I => \N__35792\
        );

    \I__6514\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35789\
        );

    \I__6513\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35774\
        );

    \I__6512\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35774\
        );

    \I__6511\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35774\
        );

    \I__6510\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35774\
        );

    \I__6509\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35774\
        );

    \I__6508\ : InMux
    port map (
            O => \N__35823\,
            I => \N__35774\
        );

    \I__6507\ : InMux
    port map (
            O => \N__35822\,
            I => \N__35774\
        );

    \I__6506\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35771\
        );

    \I__6505\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35762\
        );

    \I__6504\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35762\
        );

    \I__6503\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35762\
        );

    \I__6502\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35762\
        );

    \I__6501\ : InMux
    port map (
            O => \N__35816\,
            I => \N__35749\
        );

    \I__6500\ : InMux
    port map (
            O => \N__35815\,
            I => \N__35749\
        );

    \I__6499\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35749\
        );

    \I__6498\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35749\
        );

    \I__6497\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35749\
        );

    \I__6496\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35749\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__35806\,
            I => \N__35744\
        );

    \I__6494\ : Span4Mux_h
    port map (
            O => \N__35803\,
            I => \N__35744\
        );

    \I__6493\ : Span4Mux_v
    port map (
            O => \N__35800\,
            I => \N__35737\
        );

    \I__6492\ : Span4Mux_h
    port map (
            O => \N__35797\,
            I => \N__35737\
        );

    \I__6491\ : Span4Mux_h
    port map (
            O => \N__35792\,
            I => \N__35737\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__35789\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__35774\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__35771\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__35762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__35749\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6485\ : Odrv4
    port map (
            O => \N__35744\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6484\ : Odrv4
    port map (
            O => \N__35737\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6483\ : InMux
    port map (
            O => \N__35722\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__6482\ : IoInMux
    port map (
            O => \N__35719\,
            I => \N__35716\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__35716\,
            I => \N__35713\
        );

    \I__6480\ : Span4Mux_s0_v
    port map (
            O => \N__35713\,
            I => \N__35710\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__35710\,
            I => \GB_BUFFER_reset_c_g_THRU_CO\
        );

    \I__6478\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35701\
        );

    \I__6477\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35701\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__35701\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\
        );

    \I__6475\ : InMux
    port map (
            O => \N__35698\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__6474\ : CascadeMux
    port map (
            O => \N__35695\,
            I => \N__35692\
        );

    \I__6473\ : InMux
    port map (
            O => \N__35692\,
            I => \N__35689\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35686\
        );

    \I__6471\ : Span4Mux_h
    port map (
            O => \N__35686\,
            I => \N__35680\
        );

    \I__6470\ : InMux
    port map (
            O => \N__35685\,
            I => \N__35677\
        );

    \I__6469\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35672\
        );

    \I__6468\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35672\
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__35680\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__35677\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__35672\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__6464\ : InMux
    port map (
            O => \N__35665\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__6463\ : InMux
    port map (
            O => \N__35662\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__35659\,
            I => \N__35656\
        );

    \I__6461\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35653\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__35653\,
            I => \N__35649\
        );

    \I__6459\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35646\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__35649\,
            I => \N__35639\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__35646\,
            I => \N__35639\
        );

    \I__6456\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35636\
        );

    \I__6455\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35633\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__35639\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__35636\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__35633\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__6451\ : InMux
    port map (
            O => \N__35626\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__35623\,
            I => \N__35620\
        );

    \I__6449\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35617\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__35617\,
            I => \N__35613\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__35616\,
            I => \N__35608\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__35613\,
            I => \N__35605\
        );

    \I__6445\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35602\
        );

    \I__6444\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35597\
        );

    \I__6443\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35597\
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__35605\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__35602\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__35597\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__6439\ : InMux
    port map (
            O => \N__35590\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__6438\ : CascadeMux
    port map (
            O => \N__35587\,
            I => \N__35584\
        );

    \I__6437\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35581\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__35581\,
            I => \N__35578\
        );

    \I__6435\ : Span4Mux_h
    port map (
            O => \N__35578\,
            I => \N__35572\
        );

    \I__6434\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35569\
        );

    \I__6433\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35564\
        );

    \I__6432\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35564\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__35572\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__35569\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__35564\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__6428\ : InMux
    port map (
            O => \N__35557\,
            I => \bfn_12_23_0_\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__35554\,
            I => \N__35551\
        );

    \I__6426\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35548\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35543\
        );

    \I__6424\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35540\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__35546\,
            I => \N__35537\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__35543\,
            I => \N__35531\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__35540\,
            I => \N__35531\
        );

    \I__6420\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35526\
        );

    \I__6419\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35526\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__35531\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__35526\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__6416\ : InMux
    port map (
            O => \N__35521\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__6415\ : CascadeMux
    port map (
            O => \N__35518\,
            I => \N__35515\
        );

    \I__6414\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35511\
        );

    \I__6413\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35508\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__35511\,
            I => \N__35505\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35500\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__35505\,
            I => \N__35497\
        );

    \I__6409\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35494\
        );

    \I__6408\ : InMux
    port map (
            O => \N__35503\,
            I => \N__35491\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__35500\,
            I => \N__35488\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__35497\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__35494\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__35491\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__35488\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6402\ : InMux
    port map (
            O => \N__35479\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__35476\,
            I => \N__35473\
        );

    \I__6400\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35469\
        );

    \I__6399\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35466\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35463\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__35466\,
            I => \N__35458\
        );

    \I__6396\ : Span4Mux_h
    port map (
            O => \N__35463\,
            I => \N__35455\
        );

    \I__6395\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35452\
        );

    \I__6394\ : InMux
    port map (
            O => \N__35461\,
            I => \N__35449\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__35458\,
            I => \N__35446\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__35455\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__35452\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__35449\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__35446\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__6388\ : InMux
    port map (
            O => \N__35437\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__6387\ : InMux
    port map (
            O => \N__35434\,
            I => \N__35431\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__35431\,
            I => \N__35428\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__35428\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \N__35420\
        );

    \I__6383\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35417\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__35423\,
            I => \N__35414\
        );

    \I__6381\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35410\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__35417\,
            I => \N__35407\
        );

    \I__6379\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35404\
        );

    \I__6378\ : CascadeMux
    port map (
            O => \N__35413\,
            I => \N__35401\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35394\
        );

    \I__6376\ : Span4Mux_v
    port map (
            O => \N__35407\,
            I => \N__35394\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__35404\,
            I => \N__35394\
        );

    \I__6374\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35391\
        );

    \I__6373\ : Span4Mux_h
    port map (
            O => \N__35394\,
            I => \N__35388\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__35391\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__35388\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__6370\ : InMux
    port map (
            O => \N__35383\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__6369\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35377\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35374\
        );

    \I__6367\ : Odrv12
    port map (
            O => \N__35374\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__35371\,
            I => \N__35367\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__35370\,
            I => \N__35364\
        );

    \I__6364\ : InMux
    port map (
            O => \N__35367\,
            I => \N__35359\
        );

    \I__6363\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35356\
        );

    \I__6362\ : InMux
    port map (
            O => \N__35363\,
            I => \N__35353\
        );

    \I__6361\ : InMux
    port map (
            O => \N__35362\,
            I => \N__35350\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__35359\,
            I => \N__35345\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__35356\,
            I => \N__35345\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35342\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__35350\,
            I => \N__35339\
        );

    \I__6356\ : Span4Mux_h
    port map (
            O => \N__35345\,
            I => \N__35336\
        );

    \I__6355\ : Span4Mux_h
    port map (
            O => \N__35342\,
            I => \N__35331\
        );

    \I__6354\ : Span4Mux_h
    port map (
            O => \N__35339\,
            I => \N__35331\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__35336\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__6352\ : Odrv4
    port map (
            O => \N__35331\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__6351\ : InMux
    port map (
            O => \N__35326\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__6350\ : InMux
    port map (
            O => \N__35323\,
            I => \N__35320\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__35320\,
            I => \N__35317\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__35317\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__35314\,
            I => \N__35311\
        );

    \I__6346\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35308\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__35308\,
            I => \N__35304\
        );

    \I__6344\ : CascadeMux
    port map (
            O => \N__35307\,
            I => \N__35301\
        );

    \I__6343\ : Span4Mux_v
    port map (
            O => \N__35304\,
            I => \N__35296\
        );

    \I__6342\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35293\
        );

    \I__6341\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35290\
        );

    \I__6340\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35287\
        );

    \I__6339\ : Odrv4
    port map (
            O => \N__35296\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__35293\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__35290\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__35287\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__6335\ : InMux
    port map (
            O => \N__35278\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__6334\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35272\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__35272\,
            I => \N__35269\
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__35269\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__35266\,
            I => \N__35262\
        );

    \I__6330\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35257\
        );

    \I__6329\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35254\
        );

    \I__6328\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35251\
        );

    \I__6327\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35248\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__35257\,
            I => \N__35245\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35240\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35240\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__35248\,
            I => \N__35237\
        );

    \I__6322\ : Span4Mux_v
    port map (
            O => \N__35245\,
            I => \N__35232\
        );

    \I__6321\ : Span4Mux_h
    port map (
            O => \N__35240\,
            I => \N__35232\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__35237\,
            I => \N__35229\
        );

    \I__6319\ : Odrv4
    port map (
            O => \N__35232\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__6318\ : Odrv4
    port map (
            O => \N__35229\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__6317\ : InMux
    port map (
            O => \N__35224\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__6316\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35218\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__35218\,
            I => \N__35215\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__35215\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__35212\,
            I => \N__35209\
        );

    \I__6312\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35206\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__35206\,
            I => \N__35203\
        );

    \I__6310\ : Span4Mux_h
    port map (
            O => \N__35203\,
            I => \N__35197\
        );

    \I__6309\ : InMux
    port map (
            O => \N__35202\,
            I => \N__35194\
        );

    \I__6308\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35191\
        );

    \I__6307\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35188\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__35197\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__35194\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__35191\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__35188\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__6302\ : InMux
    port map (
            O => \N__35179\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__6301\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35173\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__35170\
        );

    \I__6299\ : Odrv4
    port map (
            O => \N__35170\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__6298\ : InMux
    port map (
            O => \N__35167\,
            I => \bfn_12_22_0_\
        );

    \I__6297\ : CascadeMux
    port map (
            O => \N__35164\,
            I => \N__35161\
        );

    \I__6296\ : InMux
    port map (
            O => \N__35161\,
            I => \N__35158\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__35158\,
            I => \N__35154\
        );

    \I__6294\ : CascadeMux
    port map (
            O => \N__35157\,
            I => \N__35151\
        );

    \I__6293\ : Span4Mux_h
    port map (
            O => \N__35154\,
            I => \N__35146\
        );

    \I__6292\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35143\
        );

    \I__6291\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35140\
        );

    \I__6290\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35137\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__35146\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__35143\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__35140\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__35137\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__6285\ : InMux
    port map (
            O => \N__35128\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__6284\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35122\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__35122\,
            I => \N__35119\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__35119\,
            I => \N__35116\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__35116\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__6280\ : InMux
    port map (
            O => \N__35113\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__6279\ : InMux
    port map (
            O => \N__35110\,
            I => \N__35107\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__35107\,
            I => \N__35104\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__35104\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__6276\ : CascadeMux
    port map (
            O => \N__35101\,
            I => \N__35098\
        );

    \I__6275\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35095\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__35095\,
            I => \N__35091\
        );

    \I__6273\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35086\
        );

    \I__6272\ : Span4Mux_h
    port map (
            O => \N__35091\,
            I => \N__35083\
        );

    \I__6271\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35080\
        );

    \I__6270\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35077\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__35086\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__35083\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__35080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__35077\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__6265\ : InMux
    port map (
            O => \N__35068\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__6264\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35062\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__35062\,
            I => \N__35059\
        );

    \I__6262\ : Odrv12
    port map (
            O => \N__35059\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__35056\,
            I => \N__35053\
        );

    \I__6260\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35048\
        );

    \I__6259\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35045\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__35051\,
            I => \N__35042\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__35038\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__35045\,
            I => \N__35035\
        );

    \I__6255\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35032\
        );

    \I__6254\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35029\
        );

    \I__6253\ : Span4Mux_h
    port map (
            O => \N__35038\,
            I => \N__35026\
        );

    \I__6252\ : Span4Mux_h
    port map (
            O => \N__35035\,
            I => \N__35023\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__35032\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__35029\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__6249\ : Odrv4
    port map (
            O => \N__35026\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__35023\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__6247\ : InMux
    port map (
            O => \N__35014\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__6246\ : InMux
    port map (
            O => \N__35011\,
            I => \N__35008\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__35008\,
            I => \N__35005\
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__35005\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__35002\,
            I => \N__34999\
        );

    \I__6242\ : InMux
    port map (
            O => \N__34999\,
            I => \N__34994\
        );

    \I__6241\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34991\
        );

    \I__6240\ : InMux
    port map (
            O => \N__34997\,
            I => \N__34987\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__34994\,
            I => \N__34984\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__34991\,
            I => \N__34981\
        );

    \I__6237\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34978\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34971\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__34984\,
            I => \N__34971\
        );

    \I__6234\ : Span4Mux_v
    port map (
            O => \N__34981\,
            I => \N__34971\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__34978\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__34971\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__6231\ : InMux
    port map (
            O => \N__34966\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__6230\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34960\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__34960\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__6228\ : CascadeMux
    port map (
            O => \N__34957\,
            I => \N__34954\
        );

    \I__6227\ : InMux
    port map (
            O => \N__34954\,
            I => \N__34951\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__34951\,
            I => \N__34947\
        );

    \I__6225\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34942\
        );

    \I__6224\ : Span4Mux_h
    port map (
            O => \N__34947\,
            I => \N__34939\
        );

    \I__6223\ : InMux
    port map (
            O => \N__34946\,
            I => \N__34936\
        );

    \I__6222\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34933\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__34942\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__34939\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__34936\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__34933\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__6217\ : InMux
    port map (
            O => \N__34924\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__6216\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34917\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__34920\,
            I => \N__34914\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__34917\,
            I => \N__34910\
        );

    \I__6213\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34906\
        );

    \I__6212\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34903\
        );

    \I__6211\ : Span4Mux_v
    port map (
            O => \N__34910\,
            I => \N__34900\
        );

    \I__6210\ : InMux
    port map (
            O => \N__34909\,
            I => \N__34897\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__34906\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__34903\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__34900\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__34897\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__34888\,
            I => \N__34885\
        );

    \I__6204\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34882\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__34882\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__6202\ : InMux
    port map (
            O => \N__34879\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__6201\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34873\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__34873\,
            I => \N__34870\
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__34870\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__34867\,
            I => \N__34864\
        );

    \I__6197\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34861\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34856\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__34860\,
            I => \N__34852\
        );

    \I__6194\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34849\
        );

    \I__6193\ : Span4Mux_h
    port map (
            O => \N__34856\,
            I => \N__34846\
        );

    \I__6192\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34843\
        );

    \I__6191\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34840\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__34849\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__34846\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__34843\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__34840\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__6186\ : InMux
    port map (
            O => \N__34831\,
            I => \bfn_12_21_0_\
        );

    \I__6185\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34825\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__34825\,
            I => \N__34819\
        );

    \I__6183\ : InMux
    port map (
            O => \N__34824\,
            I => \N__34816\
        );

    \I__6182\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34813\
        );

    \I__6181\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34810\
        );

    \I__6180\ : Span4Mux_h
    port map (
            O => \N__34819\,
            I => \N__34803\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34803\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__34813\,
            I => \N__34803\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__34810\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__6176\ : Odrv4
    port map (
            O => \N__34803\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__34798\,
            I => \N__34795\
        );

    \I__6174\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34792\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__34792\,
            I => \N__34789\
        );

    \I__6172\ : Odrv12
    port map (
            O => \N__34789\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__6171\ : InMux
    port map (
            O => \N__34786\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__6170\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34780\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__34780\,
            I => \N__34777\
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__34777\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__34774\,
            I => \N__34771\
        );

    \I__6166\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34767\
        );

    \I__6165\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34763\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__34767\,
            I => \N__34760\
        );

    \I__6163\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34756\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__34763\,
            I => \N__34753\
        );

    \I__6161\ : Span4Mux_h
    port map (
            O => \N__34760\,
            I => \N__34750\
        );

    \I__6160\ : InMux
    port map (
            O => \N__34759\,
            I => \N__34747\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__34756\,
            I => \N__34744\
        );

    \I__6158\ : Span4Mux_h
    port map (
            O => \N__34753\,
            I => \N__34741\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__34750\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__34747\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6155\ : Odrv4
    port map (
            O => \N__34744\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6154\ : Odrv4
    port map (
            O => \N__34741\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__6153\ : InMux
    port map (
            O => \N__34732\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__6152\ : InMux
    port map (
            O => \N__34729\,
            I => \N__34726\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__34726\,
            I => \N__34722\
        );

    \I__6150\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34719\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__34722\,
            I => \N__34716\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__34719\,
            I => \N__34713\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__34716\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__34713\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__34708\,
            I => \N__34705\
        );

    \I__6144\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34702\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__34702\,
            I => \N__34698\
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__34701\,
            I => \N__34694\
        );

    \I__6141\ : Span4Mux_h
    port map (
            O => \N__34698\,
            I => \N__34690\
        );

    \I__6140\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34685\
        );

    \I__6139\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34685\
        );

    \I__6138\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34682\
        );

    \I__6137\ : Odrv4
    port map (
            O => \N__34690\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__34685\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__34682\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__6134\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34672\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__34672\,
            I => \N__34669\
        );

    \I__6132\ : Odrv4
    port map (
            O => \N__34669\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__34666\,
            I => \N__34663\
        );

    \I__6130\ : InMux
    port map (
            O => \N__34663\,
            I => \N__34660\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__34660\,
            I => \N__34657\
        );

    \I__6128\ : Span4Mux_h
    port map (
            O => \N__34657\,
            I => \N__34652\
        );

    \I__6127\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34649\
        );

    \I__6126\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34646\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__34652\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__34649\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__34646\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__6122\ : InMux
    port map (
            O => \N__34639\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__6121\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34633\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__6119\ : Span4Mux_v
    port map (
            O => \N__34630\,
            I => \N__34624\
        );

    \I__6118\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34621\
        );

    \I__6117\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34618\
        );

    \I__6116\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34615\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__34624\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__34621\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__34618\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__34615\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__34606\,
            I => \N__34603\
        );

    \I__6110\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34600\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__34600\,
            I => \N__34597\
        );

    \I__6108\ : Odrv4
    port map (
            O => \N__34597\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__6107\ : InMux
    port map (
            O => \N__34594\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__6106\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34588\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__34588\,
            I => \N__34585\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__34585\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt28\
        );

    \I__6103\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34578\
        );

    \I__6102\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34575\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__34578\,
            I => \N__34572\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34569\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__34572\,
            I => \N__34566\
        );

    \I__6098\ : Span4Mux_h
    port map (
            O => \N__34569\,
            I => \N__34563\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__34566\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_28
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__34563\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_28
        );

    \I__6095\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34553\
        );

    \I__6094\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34548\
        );

    \I__6093\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34548\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__34553\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__34548\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_29\
        );

    \I__6090\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34538\
        );

    \I__6089\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34533\
        );

    \I__6088\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34533\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__34538\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_28\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__34533\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_28\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__34528\,
            I => \N__34525\
        );

    \I__6084\ : InMux
    port map (
            O => \N__34525\,
            I => \N__34522\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34522\,
            I => \N__34519\
        );

    \I__6082\ : Odrv4
    port map (
            O => \N__34519\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\
        );

    \I__6081\ : CascadeMux
    port map (
            O => \N__34516\,
            I => \N__34513\
        );

    \I__6080\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34510\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__34510\,
            I => \N__34507\
        );

    \I__6078\ : Odrv12
    port map (
            O => \N__34507\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\
        );

    \I__6077\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34499\
        );

    \I__6076\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34494\
        );

    \I__6075\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34494\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__34499\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__34494\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_30\
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__34489\,
            I => \N__34486\
        );

    \I__6071\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34474\
        );

    \I__6070\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34474\
        );

    \I__6069\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34474\
        );

    \I__6068\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34474\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__34474\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\
        );

    \I__6066\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34466\
        );

    \I__6065\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34461\
        );

    \I__6064\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34461\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__34466\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__34461\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_31\
        );

    \I__6061\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34453\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__34453\,
            I => \N__34450\
        );

    \I__6059\ : Odrv4
    port map (
            O => \N__34450\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt30\
        );

    \I__6058\ : InMux
    port map (
            O => \N__34447\,
            I => \N__34444\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__34441\,
            I => \N__34437\
        );

    \I__6055\ : InMux
    port map (
            O => \N__34440\,
            I => \N__34431\
        );

    \I__6054\ : Span4Mux_v
    port map (
            O => \N__34437\,
            I => \N__34427\
        );

    \I__6053\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34422\
        );

    \I__6052\ : InMux
    port map (
            O => \N__34435\,
            I => \N__34422\
        );

    \I__6051\ : InMux
    port map (
            O => \N__34434\,
            I => \N__34419\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__34431\,
            I => \N__34416\
        );

    \I__6049\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34413\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__34427\,
            I => \N__34410\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__34422\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__34419\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__34416\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__34413\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__34410\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6042\ : InMux
    port map (
            O => \N__34399\,
            I => \N__34392\
        );

    \I__6041\ : InMux
    port map (
            O => \N__34398\,
            I => \N__34387\
        );

    \I__6040\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34387\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__34396\,
            I => \N__34383\
        );

    \I__6038\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34380\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34377\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34374\
        );

    \I__6035\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34371\
        );

    \I__6034\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34368\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34363\
        );

    \I__6032\ : Span12Mux_h
    port map (
            O => \N__34377\,
            I => \N__34363\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__34374\,
            I => \N__34360\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__34371\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__34368\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6028\ : Odrv12
    port map (
            O => \N__34363\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__34360\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6026\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34348\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34345\
        );

    \I__6024\ : Sp12to4
    port map (
            O => \N__34345\,
            I => \N__34342\
        );

    \I__6023\ : Span12Mux_v
    port map (
            O => \N__34342\,
            I => \N__34339\
        );

    \I__6022\ : Odrv12
    port map (
            O => \N__34339\,
            I => \phase_controller_inst2.stoper_hc.un4_start_0\
        );

    \I__6021\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34330\
        );

    \I__6020\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34330\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34327\
        );

    \I__6018\ : Span4Mux_h
    port map (
            O => \N__34327\,
            I => \N__34323\
        );

    \I__6017\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34320\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__34323\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__34320\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__6014\ : InMux
    port map (
            O => \N__34315\,
            I => \N__34312\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__34312\,
            I => \N__34307\
        );

    \I__6012\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34304\
        );

    \I__6011\ : InMux
    port map (
            O => \N__34310\,
            I => \N__34301\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__34307\,
            I => \N__34298\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__34304\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__34301\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__34298\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__6006\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34288\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34285\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__34285\,
            I => \N__34282\
        );

    \I__6003\ : Span4Mux_h
    port map (
            O => \N__34282\,
            I => \N__34278\
        );

    \I__6002\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34275\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__34278\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_14
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__34275\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_14
        );

    \I__5999\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34267\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__34267\,
            I => \N__34264\
        );

    \I__5997\ : Odrv4
    port map (
            O => \N__34264\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\
        );

    \I__5996\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34258\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__34258\,
            I => \N__34255\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__34255\,
            I => \N__34251\
        );

    \I__5993\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34248\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__34251\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_12
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__34248\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_12
        );

    \I__5990\ : InMux
    port map (
            O => \N__34243\,
            I => \N__34240\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__34240\,
            I => \N__34237\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__34237\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\
        );

    \I__5987\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34231\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__34231\,
            I => \N__34228\
        );

    \I__5985\ : Span4Mux_v
    port map (
            O => \N__34228\,
            I => \N__34224\
        );

    \I__5984\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34221\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__34224\,
            I => \N__34218\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__34221\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_15
        );

    \I__5981\ : Odrv4
    port map (
            O => \N__34218\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_15
        );

    \I__5980\ : InMux
    port map (
            O => \N__34213\,
            I => \N__34210\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__34210\,
            I => \N__34207\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__34207\,
            I => \N__34204\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__34204\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\
        );

    \I__5976\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34198\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34195\
        );

    \I__5974\ : Span4Mux_h
    port map (
            O => \N__34195\,
            I => \N__34191\
        );

    \I__5973\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34188\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__34191\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_11
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__34188\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_11
        );

    \I__5970\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__34180\,
            I => \N__34177\
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__34177\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\
        );

    \I__5967\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34171\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34168\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__34168\,
            I => \N__34164\
        );

    \I__5964\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34161\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__34164\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_8
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__34161\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_8
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__34156\,
            I => \N__34153\
        );

    \I__5960\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34150\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__34150\,
            I => \N__34147\
        );

    \I__5958\ : Span4Mux_h
    port map (
            O => \N__34147\,
            I => \N__34144\
        );

    \I__5957\ : Odrv4
    port map (
            O => \N__34144\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\
        );

    \I__5956\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34138\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34134\
        );

    \I__5954\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34131\
        );

    \I__5953\ : Span4Mux_v
    port map (
            O => \N__34134\,
            I => \N__34128\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__34131\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_9
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__34128\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_9
        );

    \I__5950\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34120\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__34117\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\
        );

    \I__5947\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__34111\,
            I => \N__34108\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__34108\,
            I => \N__34104\
        );

    \I__5944\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34101\
        );

    \I__5943\ : Odrv4
    port map (
            O => \N__34104\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_10
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__34101\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_10
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__34096\,
            I => \N__34093\
        );

    \I__5940\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34090\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__34090\,
            I => \N__34087\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__34087\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\
        );

    \I__5937\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34081\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__34081\,
            I => \N__34078\
        );

    \I__5935\ : Span12Mux_v
    port map (
            O => \N__34078\,
            I => \N__34073\
        );

    \I__5934\ : InMux
    port map (
            O => \N__34077\,
            I => \N__34068\
        );

    \I__5933\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34068\
        );

    \I__5932\ : Odrv12
    port map (
            O => \N__34073\,
            I => \phase_controller_inst2.start_flagZ0\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__34068\,
            I => \phase_controller_inst2.start_flagZ0\
        );

    \I__5930\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34059\
        );

    \I__5929\ : CascadeMux
    port map (
            O => \N__34062\,
            I => \N__34056\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__34059\,
            I => \N__34052\
        );

    \I__5927\ : InMux
    port map (
            O => \N__34056\,
            I => \N__34047\
        );

    \I__5926\ : InMux
    port map (
            O => \N__34055\,
            I => \N__34047\
        );

    \I__5925\ : Span4Mux_v
    port map (
            O => \N__34052\,
            I => \N__34044\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__34047\,
            I => \N__34039\
        );

    \I__5923\ : Span4Mux_v
    port map (
            O => \N__34044\,
            I => \N__34039\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__34039\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__5921\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34029\
        );

    \I__5920\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34020\
        );

    \I__5919\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34020\
        );

    \I__5918\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34020\
        );

    \I__5917\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34020\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__34017\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__34014\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__34017\,
            I => \N__34009\
        );

    \I__5913\ : Span4Mux_v
    port map (
            O => \N__34014\,
            I => \N__34009\
        );

    \I__5912\ : Span4Mux_v
    port map (
            O => \N__34009\,
            I => \N__34005\
        );

    \I__5911\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34002\
        );

    \I__5910\ : Sp12to4
    port map (
            O => \N__34005\,
            I => \N__33997\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__34002\,
            I => \N__33997\
        );

    \I__5908\ : Span12Mux_h
    port map (
            O => \N__33997\,
            I => \N__33994\
        );

    \I__5907\ : Odrv12
    port map (
            O => \N__33994\,
            I => start_stop_c
        );

    \I__5906\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33986\
        );

    \I__5905\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33981\
        );

    \I__5904\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33981\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__33986\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__33981\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__33976\,
            I => \phase_controller_inst1.state_ns_0_0_1_cascade_\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__33973\,
            I => \N__33969\
        );

    \I__5899\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33965\
        );

    \I__5898\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33960\
        );

    \I__5897\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33960\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__33965\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__33960\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__33955\,
            I => \phase_controller_inst1.stoper_tr.un4_start_0_cascade_\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__33952\,
            I => \N__33947\
        );

    \I__5892\ : CascadeMux
    port map (
            O => \N__33951\,
            I => \N__33944\
        );

    \I__5891\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33937\
        );

    \I__5890\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33937\
        );

    \I__5889\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33937\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__33937\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__5887\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33928\
        );

    \I__5886\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33928\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__33928\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5884\ : InMux
    port map (
            O => \N__33925\,
            I => \N__33922\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__33922\,
            I => \N__33919\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__33919\,
            I => \N__33916\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__33916\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\
        );

    \I__5880\ : InMux
    port map (
            O => \N__33913\,
            I => \N__33901\
        );

    \I__5879\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33901\
        );

    \I__5878\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33901\
        );

    \I__5877\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33901\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__33901\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\
        );

    \I__5875\ : InMux
    port map (
            O => \N__33898\,
            I => \N__33893\
        );

    \I__5874\ : InMux
    port map (
            O => \N__33897\,
            I => \N__33888\
        );

    \I__5873\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33888\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__33893\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__33888\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_31\
        );

    \I__5870\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33878\
        );

    \I__5869\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33875\
        );

    \I__5868\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33872\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__33878\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__33875\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__33872\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_30\
        );

    \I__5864\ : CascadeMux
    port map (
            O => \N__33865\,
            I => \N__33862\
        );

    \I__5863\ : InMux
    port map (
            O => \N__33862\,
            I => \N__33859\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__33859\,
            I => \N__33856\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__33856\,
            I => \N__33853\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__33853\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt30\
        );

    \I__5859\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33847\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33844\
        );

    \I__5857\ : Span4Mux_h
    port map (
            O => \N__33844\,
            I => \N__33840\
        );

    \I__5856\ : InMux
    port map (
            O => \N__33843\,
            I => \N__33837\
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__33840\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__33837\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5853\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33829\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__33829\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__5851\ : CascadeMux
    port map (
            O => \N__33826\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__5850\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33820\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__33820\,
            I => \N__33817\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__33817\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\
        );

    \I__5847\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33811\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__33811\,
            I => \N__33808\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__33808\,
            I => \N__33804\
        );

    \I__5844\ : InMux
    port map (
            O => \N__33807\,
            I => \N__33801\
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__33804\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__33801\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__5841\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33793\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33789\
        );

    \I__5839\ : InMux
    port map (
            O => \N__33792\,
            I => \N__33786\
        );

    \I__5838\ : Span12Mux_v
    port map (
            O => \N__33789\,
            I => \N__33783\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__33786\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__5836\ : Odrv12
    port map (
            O => \N__33783\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__5835\ : InMux
    port map (
            O => \N__33778\,
            I => \N__33773\
        );

    \I__5834\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33762\
        );

    \I__5833\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33762\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__33773\,
            I => \N__33759\
        );

    \I__5831\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33754\
        );

    \I__5830\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33754\
        );

    \I__5829\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33744\
        );

    \I__5828\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33744\
        );

    \I__5827\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33741\
        );

    \I__5826\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33738\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33735\
        );

    \I__5824\ : Span4Mux_h
    port map (
            O => \N__33759\,
            I => \N__33730\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__33754\,
            I => \N__33730\
        );

    \I__5822\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33714\
        );

    \I__5821\ : InMux
    port map (
            O => \N__33752\,
            I => \N__33714\
        );

    \I__5820\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33714\
        );

    \I__5819\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33714\
        );

    \I__5818\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33711\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33704\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33704\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33699\
        );

    \I__5814\ : Span4Mux_v
    port map (
            O => \N__33735\,
            I => \N__33699\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__33730\,
            I => \N__33696\
        );

    \I__5812\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33686\
        );

    \I__5811\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33686\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__33727\,
            I => \N__33683\
        );

    \I__5809\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33672\
        );

    \I__5808\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33672\
        );

    \I__5807\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33672\
        );

    \I__5806\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33672\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__33714\,
            I => \N__33667\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__33711\,
            I => \N__33667\
        );

    \I__5803\ : InMux
    port map (
            O => \N__33710\,
            I => \N__33662\
        );

    \I__5802\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33662\
        );

    \I__5801\ : Span4Mux_v
    port map (
            O => \N__33704\,
            I => \N__33659\
        );

    \I__5800\ : Sp12to4
    port map (
            O => \N__33699\,
            I => \N__33654\
        );

    \I__5799\ : Sp12to4
    port map (
            O => \N__33696\,
            I => \N__33654\
        );

    \I__5798\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33649\
        );

    \I__5797\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33649\
        );

    \I__5796\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33642\
        );

    \I__5795\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33642\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33642\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__33686\,
            I => \N__33639\
        );

    \I__5792\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33632\
        );

    \I__5791\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33632\
        );

    \I__5790\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33632\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33627\
        );

    \I__5788\ : Span4Mux_h
    port map (
            O => \N__33667\,
            I => \N__33627\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33662\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5786\ : Odrv4
    port map (
            O => \N__33659\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5785\ : Odrv12
    port map (
            O => \N__33654\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__33649\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__33642\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5782\ : Odrv12
    port map (
            O => \N__33639\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__33632\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__33627\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__5779\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33604\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__33604\,
            I => \N__33600\
        );

    \I__5776\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33597\
        );

    \I__5775\ : Odrv4
    port map (
            O => \N__33600\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__33597\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__5773\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33589\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__33589\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__33586\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\
        );

    \I__5770\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33580\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__5768\ : Span4Mux_h
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__33574\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\
        );

    \I__5766\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33565\
        );

    \I__5765\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33565\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__33565\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\
        );

    \I__5763\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33555\
        );

    \I__5762\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33555\
        );

    \I__5761\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33552\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__33555\,
            I => \N__33549\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__33552\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_25\
        );

    \I__5758\ : Odrv4
    port map (
            O => \N__33549\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_25\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__33544\,
            I => \N__33540\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__33543\,
            I => \N__33537\
        );

    \I__5755\ : InMux
    port map (
            O => \N__33540\,
            I => \N__33532\
        );

    \I__5754\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33532\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__33532\,
            I => \N__33529\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__33529\,
            I => \N__33526\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__33526\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\
        );

    \I__5750\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33516\
        );

    \I__5749\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33516\
        );

    \I__5748\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33513\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__33516\,
            I => \N__33510\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__33513\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_24\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__33510\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_24\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__33505\,
            I => \N__33502\
        );

    \I__5743\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__33499\,
            I => \N__33496\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__33496\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\
        );

    \I__5740\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33490\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__33490\,
            I => \N__33487\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__33487\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt26\
        );

    \I__5737\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33478\
        );

    \I__5736\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33478\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__33478\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\
        );

    \I__5734\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33468\
        );

    \I__5733\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33468\
        );

    \I__5732\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33465\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__33468\,
            I => \N__33462\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__33465\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_27\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__33462\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_27\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__33457\,
            I => \N__33453\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__33456\,
            I => \N__33450\
        );

    \I__5726\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33445\
        );

    \I__5725\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33445\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__33445\,
            I => \N__33441\
        );

    \I__5723\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33438\
        );

    \I__5722\ : Span4Mux_v
    port map (
            O => \N__33441\,
            I => \N__33435\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__33438\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_26\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__33435\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_26\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__33430\,
            I => \N__33427\
        );

    \I__5718\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33424\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__33424\,
            I => \N__33421\
        );

    \I__5716\ : Span4Mux_h
    port map (
            O => \N__33421\,
            I => \N__33418\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__33418\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\
        );

    \I__5714\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33409\
        );

    \I__5713\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33409\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__33409\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\
        );

    \I__5711\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33403\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__33403\,
            I => \N__33400\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__33400\,
            I => \N__33397\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__33397\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt28\
        );

    \I__5707\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33389\
        );

    \I__5706\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33384\
        );

    \I__5705\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33384\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__33389\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_29\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__33384\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_29\
        );

    \I__5702\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33374\
        );

    \I__5701\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33369\
        );

    \I__5700\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33369\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__33374\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_28\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__33369\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_28\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__33364\,
            I => \N__33361\
        );

    \I__5696\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33358\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__33358\,
            I => \N__33355\
        );

    \I__5694\ : Span4Mux_v
    port map (
            O => \N__33355\,
            I => \N__33352\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__33352\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\
        );

    \I__5692\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33343\
        );

    \I__5691\ : InMux
    port map (
            O => \N__33348\,
            I => \N__33343\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__33343\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\
        );

    \I__5689\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33334\
        );

    \I__5688\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33334\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__33334\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\
        );

    \I__5686\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33325\
        );

    \I__5685\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33325\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__33325\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\
        );

    \I__5683\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33310\
        );

    \I__5682\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33310\
        );

    \I__5681\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33310\
        );

    \I__5680\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33310\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__33310\,
            I => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\
        );

    \I__5678\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33304\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__33304\,
            I => \N__33301\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__33301\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt24\
        );

    \I__5675\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33295\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__33295\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\
        );

    \I__5673\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33289\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__33289\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\
        );

    \I__5671\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33283\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__33283\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt16\
        );

    \I__5669\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33274\
        );

    \I__5668\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33274\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__33274\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\
        );

    \I__5666\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33265\
        );

    \I__5665\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33265\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__33265\,
            I => \N__33261\
        );

    \I__5663\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33258\
        );

    \I__5662\ : Span4Mux_h
    port map (
            O => \N__33261\,
            I => \N__33255\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__33258\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_17\
        );

    \I__5660\ : Odrv4
    port map (
            O => \N__33255\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_17\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__33250\,
            I => \N__33246\
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__33249\,
            I => \N__33243\
        );

    \I__5657\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33238\
        );

    \I__5656\ : InMux
    port map (
            O => \N__33243\,
            I => \N__33238\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33234\
        );

    \I__5654\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33231\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__33234\,
            I => \N__33228\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__33231\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_16\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__33228\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_16\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__33223\,
            I => \N__33220\
        );

    \I__5649\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33217\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__33217\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\
        );

    \I__5647\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33208\
        );

    \I__5646\ : InMux
    port map (
            O => \N__33213\,
            I => \N__33208\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__33208\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\
        );

    \I__5644\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33201\
        );

    \I__5643\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33198\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33195\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__33198\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__33195\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\
        );

    \I__5639\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33186\
        );

    \I__5638\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33182\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33179\
        );

    \I__5636\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33176\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__33182\,
            I => \N__33171\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__33179\,
            I => \N__33171\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__33176\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__33171\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_19\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__33166\,
            I => \N__33162\
        );

    \I__5630\ : CascadeMux
    port map (
            O => \N__33165\,
            I => \N__33159\
        );

    \I__5629\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33156\
        );

    \I__5628\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33153\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33149\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__33153\,
            I => \N__33146\
        );

    \I__5625\ : InMux
    port map (
            O => \N__33152\,
            I => \N__33143\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__33149\,
            I => \N__33140\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__33146\,
            I => \N__33137\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__33143\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__33140\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__33137\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_18\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__33130\,
            I => \N__33127\
        );

    \I__5618\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33124\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__33124\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\
        );

    \I__5616\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33117\
        );

    \I__5615\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33114\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__33117\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__33114\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\
        );

    \I__5612\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33103\
        );

    \I__5611\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33103\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__33103\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\
        );

    \I__5609\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__33097\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\
        );

    \I__5607\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__33091\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\
        );

    \I__5605\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33085\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__33085\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\
        );

    \I__5603\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__33079\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__33076\,
            I => \N__33073\
        );

    \I__5600\ : InMux
    port map (
            O => \N__33073\,
            I => \N__33070\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__33070\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\
        );

    \I__5598\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33064\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__33064\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\
        );

    \I__5596\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33058\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__33058\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\
        );

    \I__5594\ : InMux
    port map (
            O => \N__33055\,
            I => \N__33052\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__33052\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\
        );

    \I__5592\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33046\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__33046\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__33043\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\
        );

    \I__5589\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33037\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__33037\,
            I => \N__33034\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__33034\,
            I => \current_shift_inst.PI_CTRL.N_46_21\
        );

    \I__5586\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__33025\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__33025\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__5583\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33019\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__33019\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__5581\ : InMux
    port map (
            O => \N__33016\,
            I => \N__33013\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__33013\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__5579\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__33007\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\
        );

    \I__5577\ : InMux
    port map (
            O => \N__33004\,
            I => \N__33001\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__33001\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\
        );

    \I__5575\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__32995\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\
        );

    \I__5573\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32989\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__32989\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__32986\,
            I => \N__32983\
        );

    \I__5570\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32980\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__32980\,
            I => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\
        );

    \I__5568\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__32968\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__32965\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\
        );

    \I__5563\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32959\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__32959\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__32956\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\
        );

    \I__5560\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32950\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__32950\,
            I => \current_shift_inst.PI_CTRL.N_77\
        );

    \I__5558\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__32944\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__32941\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\
        );

    \I__5555\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32935\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__32935\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\
        );

    \I__5553\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32929\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__32929\,
            I => \current_shift_inst.PI_CTRL.N_46_16\
        );

    \I__5551\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32919\
        );

    \I__5550\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32919\
        );

    \I__5549\ : CEMux
    port map (
            O => \N__32924\,
            I => \N__32895\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32892\
        );

    \I__5547\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32883\
        );

    \I__5546\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32883\
        );

    \I__5545\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32883\
        );

    \I__5544\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32883\
        );

    \I__5543\ : InMux
    port map (
            O => \N__32914\,
            I => \N__32874\
        );

    \I__5542\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32871\
        );

    \I__5541\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32858\
        );

    \I__5540\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32858\
        );

    \I__5539\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32858\
        );

    \I__5538\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32858\
        );

    \I__5537\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32858\
        );

    \I__5536\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32858\
        );

    \I__5535\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32843\
        );

    \I__5534\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32843\
        );

    \I__5533\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32843\
        );

    \I__5532\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32843\
        );

    \I__5531\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32843\
        );

    \I__5530\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32843\
        );

    \I__5529\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32843\
        );

    \I__5528\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32838\
        );

    \I__5527\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32838\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32835\
        );

    \I__5525\ : Span4Mux_v
    port map (
            O => \N__32892\,
            I => \N__32830\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32830\
        );

    \I__5523\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32825\
        );

    \I__5522\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32825\
        );

    \I__5521\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32822\
        );

    \I__5520\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32819\
        );

    \I__5519\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32814\
        );

    \I__5518\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32814\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__32874\,
            I => \N__32811\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32808\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__32858\,
            I => \N__32803\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32803\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__32838\,
            I => \N__32796\
        );

    \I__5512\ : Span4Mux_v
    port map (
            O => \N__32835\,
            I => \N__32796\
        );

    \I__5511\ : Span4Mux_v
    port map (
            O => \N__32830\,
            I => \N__32796\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__32825\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__32822\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__32819\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__32814\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5506\ : Odrv12
    port map (
            O => \N__32811\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5505\ : Odrv4
    port map (
            O => \N__32808\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__32803\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__32796\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__5502\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32776\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__32776\,
            I => \N__32773\
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__32773\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__32770\,
            I => \N__32767\
        );

    \I__5498\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32764\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__32764\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt22\
        );

    \I__5496\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32758\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__32758\,
            I => \N__32755\
        );

    \I__5494\ : Span4Mux_h
    port map (
            O => \N__32755\,
            I => \N__32751\
        );

    \I__5493\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32748\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__32751\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_22
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__32748\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_22
        );

    \I__5490\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32736\
        );

    \I__5489\ : InMux
    port map (
            O => \N__32742\,
            I => \N__32736\
        );

    \I__5488\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32733\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__32736\,
            I => \N__32730\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__32733\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__32730\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_23\
        );

    \I__5484\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32719\
        );

    \I__5483\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32719\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__32719\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\
        );

    \I__5481\ : CascadeMux
    port map (
            O => \N__32716\,
            I => \N__32712\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__32715\,
            I => \N__32709\
        );

    \I__5479\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32703\
        );

    \I__5478\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32703\
        );

    \I__5477\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32700\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32697\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__32700\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__32697\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_22\
        );

    \I__5473\ : InMux
    port map (
            O => \N__32692\,
            I => \N__32689\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__32689\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\
        );

    \I__5471\ : InMux
    port map (
            O => \N__32686\,
            I => \N__32683\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__32683\,
            I => \N__32680\
        );

    \I__5469\ : Span4Mux_h
    port map (
            O => \N__32680\,
            I => \N__32676\
        );

    \I__5468\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32673\
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__32676\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_23
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__32673\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_23
        );

    \I__5465\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32662\
        );

    \I__5464\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32662\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__32662\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\
        );

    \I__5462\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32647\
        );

    \I__5461\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32647\
        );

    \I__5460\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32647\
        );

    \I__5459\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32647\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32644\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__32644\,
            I => \N__32641\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__32641\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\
        );

    \I__5455\ : CEMux
    port map (
            O => \N__32638\,
            I => \N__32632\
        );

    \I__5454\ : CEMux
    port map (
            O => \N__32637\,
            I => \N__32629\
        );

    \I__5453\ : CEMux
    port map (
            O => \N__32636\,
            I => \N__32626\
        );

    \I__5452\ : CEMux
    port map (
            O => \N__32635\,
            I => \N__32623\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32620\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__32629\,
            I => \N__32616\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32612\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32609\
        );

    \I__5447\ : Span4Mux_v
    port map (
            O => \N__32620\,
            I => \N__32606\
        );

    \I__5446\ : CEMux
    port map (
            O => \N__32619\,
            I => \N__32603\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__32616\,
            I => \N__32600\
        );

    \I__5444\ : CEMux
    port map (
            O => \N__32615\,
            I => \N__32597\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__32612\,
            I => \N__32593\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__32609\,
            I => \N__32582\
        );

    \I__5441\ : Span4Mux_h
    port map (
            O => \N__32606\,
            I => \N__32582\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32582\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__32600\,
            I => \N__32582\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__32597\,
            I => \N__32582\
        );

    \I__5437\ : CEMux
    port map (
            O => \N__32596\,
            I => \N__32579\
        );

    \I__5436\ : Span4Mux_v
    port map (
            O => \N__32593\,
            I => \N__32576\
        );

    \I__5435\ : Span4Mux_v
    port map (
            O => \N__32582\,
            I => \N__32571\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__32579\,
            I => \N__32571\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__32576\,
            I => \N__32568\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__32571\,
            I => \N__32565\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__32568\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__32565\,
            I => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\
        );

    \I__5429\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32557\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__32557\,
            I => \N__32552\
        );

    \I__5427\ : InMux
    port map (
            O => \N__32556\,
            I => \N__32549\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__32555\,
            I => \N__32546\
        );

    \I__5425\ : Span4Mux_v
    port map (
            O => \N__32552\,
            I => \N__32541\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32538\
        );

    \I__5423\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32530\
        );

    \I__5422\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32530\
        );

    \I__5421\ : InMux
    port map (
            O => \N__32544\,
            I => \N__32530\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__32541\,
            I => \N__32525\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__32538\,
            I => \N__32525\
        );

    \I__5418\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32522\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__32530\,
            I => \N__32519\
        );

    \I__5416\ : Sp12to4
    port map (
            O => \N__32525\,
            I => \N__32516\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__32522\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__32519\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__5413\ : Odrv12
    port map (
            O => \N__32516\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__5412\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32471\
        );

    \I__5411\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32471\
        );

    \I__5410\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32471\
        );

    \I__5409\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32462\
        );

    \I__5408\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32462\
        );

    \I__5407\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32462\
        );

    \I__5406\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32462\
        );

    \I__5405\ : InMux
    port map (
            O => \N__32502\,
            I => \N__32453\
        );

    \I__5404\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32453\
        );

    \I__5403\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32453\
        );

    \I__5402\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32453\
        );

    \I__5401\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32442\
        );

    \I__5400\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32442\
        );

    \I__5399\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32442\
        );

    \I__5398\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32442\
        );

    \I__5397\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32442\
        );

    \I__5396\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32433\
        );

    \I__5395\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32433\
        );

    \I__5394\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32433\
        );

    \I__5393\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32433\
        );

    \I__5392\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32424\
        );

    \I__5391\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32424\
        );

    \I__5390\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32424\
        );

    \I__5389\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32424\
        );

    \I__5388\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32415\
        );

    \I__5387\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32415\
        );

    \I__5386\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32415\
        );

    \I__5385\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32415\
        );

    \I__5384\ : InMux
    port map (
            O => \N__32481\,
            I => \N__32406\
        );

    \I__5383\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32406\
        );

    \I__5382\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32406\
        );

    \I__5381\ : InMux
    port map (
            O => \N__32478\,
            I => \N__32406\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__32471\,
            I => \N__32403\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__32462\,
            I => \N__32398\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__32453\,
            I => \N__32398\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__32442\,
            I => \N__32395\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__32433\,
            I => \N__32390\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32390\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32381\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__32406\,
            I => \N__32381\
        );

    \I__5372\ : Span4Mux_v
    port map (
            O => \N__32403\,
            I => \N__32381\
        );

    \I__5371\ : Span4Mux_v
    port map (
            O => \N__32398\,
            I => \N__32381\
        );

    \I__5370\ : Span4Mux_v
    port map (
            O => \N__32395\,
            I => \N__32374\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__32390\,
            I => \N__32374\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__32381\,
            I => \N__32374\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__32374\,
            I => \phase_controller_inst2.stoper_tr.start_latched_i_0\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__32371\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\
        );

    \I__5365\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32362\
        );

    \I__5364\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32362\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__32362\,
            I => \N__32358\
        );

    \I__5362\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32355\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__32358\,
            I => \N__32352\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__32355\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__5359\ : Odrv4
    port map (
            O => \N__32352\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_27\
        );

    \I__5358\ : InMux
    port map (
            O => \N__32347\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_26\
        );

    \I__5357\ : InMux
    port map (
            O => \N__32344\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_27\
        );

    \I__5356\ : InMux
    port map (
            O => \N__32341\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_28\
        );

    \I__5355\ : InMux
    port map (
            O => \N__32338\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_29\
        );

    \I__5354\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32303\
        );

    \I__5353\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32303\
        );

    \I__5352\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32303\
        );

    \I__5351\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32303\
        );

    \I__5350\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32294\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32294\
        );

    \I__5348\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32294\
        );

    \I__5347\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32294\
        );

    \I__5346\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32285\
        );

    \I__5345\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32285\
        );

    \I__5344\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32285\
        );

    \I__5343\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32285\
        );

    \I__5342\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32276\
        );

    \I__5341\ : InMux
    port map (
            O => \N__32322\,
            I => \N__32276\
        );

    \I__5340\ : InMux
    port map (
            O => \N__32321\,
            I => \N__32276\
        );

    \I__5339\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32276\
        );

    \I__5338\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32259\
        );

    \I__5337\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32259\
        );

    \I__5336\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32259\
        );

    \I__5335\ : InMux
    port map (
            O => \N__32316\,
            I => \N__32259\
        );

    \I__5334\ : InMux
    port map (
            O => \N__32315\,
            I => \N__32250\
        );

    \I__5333\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32250\
        );

    \I__5332\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32250\
        );

    \I__5331\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32250\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__32303\,
            I => \N__32247\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__32294\,
            I => \N__32244\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__32285\,
            I => \N__32241\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32238\
        );

    \I__5326\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32229\
        );

    \I__5325\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32229\
        );

    \I__5324\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32229\
        );

    \I__5323\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32229\
        );

    \I__5322\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32220\
        );

    \I__5321\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32220\
        );

    \I__5320\ : InMux
    port map (
            O => \N__32269\,
            I => \N__32220\
        );

    \I__5319\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32220\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__32259\,
            I => \N__32215\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__32250\,
            I => \N__32215\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__32247\,
            I => \N__32210\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__32244\,
            I => \N__32210\
        );

    \I__5314\ : Span4Mux_h
    port map (
            O => \N__32241\,
            I => \N__32205\
        );

    \I__5313\ : Span4Mux_h
    port map (
            O => \N__32238\,
            I => \N__32205\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__32229\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__32220\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__32215\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__32210\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__32205\,
            I => \phase_controller_inst1.stoper_tr.start_latched_i_0\
        );

    \I__5307\ : InMux
    port map (
            O => \N__32194\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_30\
        );

    \I__5306\ : CEMux
    port map (
            O => \N__32191\,
            I => \N__32179\
        );

    \I__5305\ : CEMux
    port map (
            O => \N__32190\,
            I => \N__32179\
        );

    \I__5304\ : CEMux
    port map (
            O => \N__32189\,
            I => \N__32179\
        );

    \I__5303\ : CEMux
    port map (
            O => \N__32188\,
            I => \N__32179\
        );

    \I__5302\ : GlobalMux
    port map (
            O => \N__32179\,
            I => \N__32176\
        );

    \I__5301\ : gio2CtrlBuf
    port map (
            O => \N__32176\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0_g\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__32173\,
            I => \N__32170\
        );

    \I__5299\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32167\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__32167\,
            I => \N__32164\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__32164\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt20\
        );

    \I__5296\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32158\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__32158\,
            I => \N__32155\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__32155\,
            I => \N__32151\
        );

    \I__5293\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32148\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__32151\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_20
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__32148\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_20
        );

    \I__5290\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32137\
        );

    \I__5289\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32137\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__32137\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\
        );

    \I__5287\ : InMux
    port map (
            O => \N__32134\,
            I => \N__32128\
        );

    \I__5286\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32128\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__32128\,
            I => \N__32125\
        );

    \I__5284\ : Odrv12
    port map (
            O => \N__32125\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__32122\,
            I => \N__32118\
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__32121\,
            I => \N__32115\
        );

    \I__5281\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32109\
        );

    \I__5280\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32109\
        );

    \I__5279\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32106\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__32109\,
            I => \N__32103\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__32106\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__32103\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_21\
        );

    \I__5275\ : InMux
    port map (
            O => \N__32098\,
            I => \N__32091\
        );

    \I__5274\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32091\
        );

    \I__5273\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32088\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32085\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__32088\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__32085\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_20\
        );

    \I__5269\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32077\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__32077\,
            I => \N__32074\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__32074\,
            I => \N__32071\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__32071\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\
        );

    \I__5265\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32061\
        );

    \I__5264\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32061\
        );

    \I__5263\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32058\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32055\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__32058\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_18\
        );

    \I__5260\ : Odrv12
    port map (
            O => \N__32055\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_18\
        );

    \I__5259\ : InMux
    port map (
            O => \N__32050\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_17\
        );

    \I__5258\ : InMux
    port map (
            O => \N__32047\,
            I => \N__32040\
        );

    \I__5257\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32040\
        );

    \I__5256\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32037\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32034\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__32037\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_19\
        );

    \I__5253\ : Odrv12
    port map (
            O => \N__32034\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_19\
        );

    \I__5252\ : InMux
    port map (
            O => \N__32029\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_18\
        );

    \I__5251\ : InMux
    port map (
            O => \N__32026\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_19\
        );

    \I__5250\ : InMux
    port map (
            O => \N__32023\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_20\
        );

    \I__5249\ : InMux
    port map (
            O => \N__32020\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_21\
        );

    \I__5248\ : InMux
    port map (
            O => \N__32017\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_22\
        );

    \I__5247\ : InMux
    port map (
            O => \N__32014\,
            I => \N__32008\
        );

    \I__5246\ : InMux
    port map (
            O => \N__32013\,
            I => \N__32008\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__32008\,
            I => \N__32004\
        );

    \I__5244\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32001\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__32004\,
            I => \N__31998\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__32001\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__5241\ : Odrv4
    port map (
            O => \N__31998\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_24\
        );

    \I__5240\ : InMux
    port map (
            O => \N__31993\,
            I => \bfn_11_16_0_\
        );

    \I__5239\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31984\
        );

    \I__5238\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31984\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__31984\,
            I => \N__31980\
        );

    \I__5236\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31977\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__31980\,
            I => \N__31974\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__31977\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__31974\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_25\
        );

    \I__5232\ : InMux
    port map (
            O => \N__31969\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_24\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__31966\,
            I => \N__31962\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__31965\,
            I => \N__31959\
        );

    \I__5229\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31954\
        );

    \I__5228\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31954\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31950\
        );

    \I__5226\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31947\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__31950\,
            I => \N__31944\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__31947\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_26\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__31944\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_26\
        );

    \I__5222\ : InMux
    port map (
            O => \N__31939\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_25\
        );

    \I__5221\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31933\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__31933\,
            I => \N__31929\
        );

    \I__5219\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31926\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__31929\,
            I => \N__31923\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__31926\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_10\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__31923\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_10\
        );

    \I__5215\ : InMux
    port map (
            O => \N__31918\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_9\
        );

    \I__5214\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31911\
        );

    \I__5213\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31908\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__31911\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_11\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__31908\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_11\
        );

    \I__5210\ : InMux
    port map (
            O => \N__31903\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_10\
        );

    \I__5209\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31896\
        );

    \I__5208\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31893\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__31896\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_12\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__31893\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_12\
        );

    \I__5205\ : InMux
    port map (
            O => \N__31888\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_11\
        );

    \I__5204\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31881\
        );

    \I__5203\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31878\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__31881\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_13\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__31878\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_13\
        );

    \I__5200\ : InMux
    port map (
            O => \N__31873\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_12\
        );

    \I__5199\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31866\
        );

    \I__5198\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31863\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__31866\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_14\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__31863\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_14\
        );

    \I__5195\ : InMux
    port map (
            O => \N__31858\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_13\
        );

    \I__5194\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31851\
        );

    \I__5193\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31848\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__31851\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_15\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__31848\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_15\
        );

    \I__5190\ : InMux
    port map (
            O => \N__31843\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_14\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__31840\,
            I => \N__31836\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__31839\,
            I => \N__31833\
        );

    \I__5187\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31828\
        );

    \I__5186\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31828\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__31828\,
            I => \N__31824\
        );

    \I__5184\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31821\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__31824\,
            I => \N__31818\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__31821\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__31818\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_16\
        );

    \I__5180\ : InMux
    port map (
            O => \N__31813\,
            I => \bfn_11_15_0_\
        );

    \I__5179\ : InMux
    port map (
            O => \N__31810\,
            I => \N__31804\
        );

    \I__5178\ : InMux
    port map (
            O => \N__31809\,
            I => \N__31804\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31800\
        );

    \I__5176\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31797\
        );

    \I__5175\ : Span4Mux_h
    port map (
            O => \N__31800\,
            I => \N__31794\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__31797\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__31794\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_17\
        );

    \I__5172\ : InMux
    port map (
            O => \N__31789\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_16\
        );

    \I__5171\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31782\
        );

    \I__5170\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31779\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__31782\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_1\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__31779\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_1\
        );

    \I__5167\ : InMux
    port map (
            O => \N__31774\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_0\
        );

    \I__5166\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31767\
        );

    \I__5165\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31764\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__31767\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_2\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__31764\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_2\
        );

    \I__5162\ : InMux
    port map (
            O => \N__31759\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_1\
        );

    \I__5161\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31752\
        );

    \I__5160\ : InMux
    port map (
            O => \N__31755\,
            I => \N__31749\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__31752\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_3\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__31749\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_3\
        );

    \I__5157\ : InMux
    port map (
            O => \N__31744\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_2\
        );

    \I__5156\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31737\
        );

    \I__5155\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31734\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__31737\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_4\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__31734\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_4\
        );

    \I__5152\ : InMux
    port map (
            O => \N__31729\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_3\
        );

    \I__5151\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31722\
        );

    \I__5150\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31719\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31716\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__31719\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_5\
        );

    \I__5147\ : Odrv4
    port map (
            O => \N__31716\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_5\
        );

    \I__5146\ : InMux
    port map (
            O => \N__31711\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_4\
        );

    \I__5145\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31704\
        );

    \I__5144\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31701\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__31704\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_6\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__31701\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_6\
        );

    \I__5141\ : InMux
    port map (
            O => \N__31696\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_5\
        );

    \I__5140\ : InMux
    port map (
            O => \N__31693\,
            I => \N__31689\
        );

    \I__5139\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31686\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__31689\,
            I => \N__31683\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__31686\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_7\
        );

    \I__5136\ : Odrv4
    port map (
            O => \N__31683\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_7\
        );

    \I__5135\ : InMux
    port map (
            O => \N__31678\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_6\
        );

    \I__5134\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31671\
        );

    \I__5133\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31668\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__31671\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_8\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__31668\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_8\
        );

    \I__5130\ : InMux
    port map (
            O => \N__31663\,
            I => \bfn_11_14_0_\
        );

    \I__5129\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31656\
        );

    \I__5128\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31653\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__31656\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_9\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__31653\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_9\
        );

    \I__5125\ : InMux
    port map (
            O => \N__31648\,
            I => \phase_controller_inst1.stoper_tr.counter_cry_8\
        );

    \I__5124\ : InMux
    port map (
            O => \N__31645\,
            I => \bfn_11_12_0_\
        );

    \I__5123\ : InMux
    port map (
            O => \N__31642\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_24\
        );

    \I__5122\ : InMux
    port map (
            O => \N__31639\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_25\
        );

    \I__5121\ : InMux
    port map (
            O => \N__31636\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_26\
        );

    \I__5120\ : InMux
    port map (
            O => \N__31633\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_27\
        );

    \I__5119\ : InMux
    port map (
            O => \N__31630\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_28\
        );

    \I__5118\ : InMux
    port map (
            O => \N__31627\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_29\
        );

    \I__5117\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31590\
        );

    \I__5116\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31590\
        );

    \I__5115\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31590\
        );

    \I__5114\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31579\
        );

    \I__5113\ : InMux
    port map (
            O => \N__31620\,
            I => \N__31579\
        );

    \I__5112\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31579\
        );

    \I__5111\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31579\
        );

    \I__5110\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31579\
        );

    \I__5109\ : InMux
    port map (
            O => \N__31616\,
            I => \N__31566\
        );

    \I__5108\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31566\
        );

    \I__5107\ : InMux
    port map (
            O => \N__31614\,
            I => \N__31566\
        );

    \I__5106\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31566\
        );

    \I__5105\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31557\
        );

    \I__5104\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31557\
        );

    \I__5103\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31557\
        );

    \I__5102\ : InMux
    port map (
            O => \N__31609\,
            I => \N__31557\
        );

    \I__5101\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31548\
        );

    \I__5100\ : InMux
    port map (
            O => \N__31607\,
            I => \N__31548\
        );

    \I__5099\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31548\
        );

    \I__5098\ : InMux
    port map (
            O => \N__31605\,
            I => \N__31548\
        );

    \I__5097\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31539\
        );

    \I__5096\ : InMux
    port map (
            O => \N__31603\,
            I => \N__31539\
        );

    \I__5095\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31539\
        );

    \I__5094\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31539\
        );

    \I__5093\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31530\
        );

    \I__5092\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31530\
        );

    \I__5091\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31530\
        );

    \I__5090\ : InMux
    port map (
            O => \N__31597\,
            I => \N__31530\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__31590\,
            I => \N__31527\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__31579\,
            I => \N__31524\
        );

    \I__5087\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31515\
        );

    \I__5086\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31515\
        );

    \I__5085\ : InMux
    port map (
            O => \N__31576\,
            I => \N__31515\
        );

    \I__5084\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31515\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31500\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__31557\,
            I => \N__31500\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__31548\,
            I => \N__31500\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__31539\,
            I => \N__31500\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31500\
        );

    \I__5078\ : Span4Mux_v
    port map (
            O => \N__31527\,
            I => \N__31500\
        );

    \I__5077\ : Span4Mux_v
    port map (
            O => \N__31524\,
            I => \N__31500\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__31515\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__31500\,
            I => \phase_controller_inst2.stoper_hc.start_latched_i_0\
        );

    \I__5074\ : InMux
    port map (
            O => \N__31495\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_30\
        );

    \I__5073\ : CEMux
    port map (
            O => \N__31492\,
            I => \N__31486\
        );

    \I__5072\ : CEMux
    port map (
            O => \N__31491\,
            I => \N__31483\
        );

    \I__5071\ : CEMux
    port map (
            O => \N__31490\,
            I => \N__31480\
        );

    \I__5070\ : CEMux
    port map (
            O => \N__31489\,
            I => \N__31477\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__31486\,
            I => \N__31474\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31469\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__31480\,
            I => \N__31469\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__31477\,
            I => \N__31466\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__31474\,
            I => \N__31463\
        );

    \I__5064\ : Span4Mux_v
    port map (
            O => \N__31469\,
            I => \N__31460\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__31466\,
            I => \N__31457\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__31463\,
            I => \N__31452\
        );

    \I__5061\ : Span4Mux_h
    port map (
            O => \N__31460\,
            I => \N__31452\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__31457\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__31452\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__31447\,
            I => \N__31443\
        );

    \I__5057\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31440\
        );

    \I__5056\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31437\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__31440\,
            I => \N__31432\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31432\
        );

    \I__5053\ : Span4Mux_v
    port map (
            O => \N__31432\,
            I => \N__31429\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__31429\,
            I => \phase_controller_inst1.stoper_tr.counter\
        );

    \I__5051\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31422\
        );

    \I__5050\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31419\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__31422\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_0\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__31419\,
            I => \phase_controller_inst1.stoper_tr.counterZ0Z_0\
        );

    \I__5047\ : InMux
    port map (
            O => \N__31414\,
            I => \bfn_11_11_0_\
        );

    \I__5046\ : InMux
    port map (
            O => \N__31411\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_16\
        );

    \I__5045\ : InMux
    port map (
            O => \N__31408\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_17\
        );

    \I__5044\ : InMux
    port map (
            O => \N__31405\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_18\
        );

    \I__5043\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31395\
        );

    \I__5042\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31395\
        );

    \I__5041\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31392\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__31395\,
            I => \N__31389\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__31392\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_20\
        );

    \I__5038\ : Odrv4
    port map (
            O => \N__31389\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_20\
        );

    \I__5037\ : InMux
    port map (
            O => \N__31384\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_19\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__31381\,
            I => \N__31377\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__31380\,
            I => \N__31374\
        );

    \I__5034\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31368\
        );

    \I__5033\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31368\
        );

    \I__5032\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31365\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__31368\,
            I => \N__31362\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__31365\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_21\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__31362\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_21\
        );

    \I__5028\ : InMux
    port map (
            O => \N__31357\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_20\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__31354\,
            I => \N__31350\
        );

    \I__5026\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31345\
        );

    \I__5025\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31345\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__31345\,
            I => \N__31341\
        );

    \I__5023\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31338\
        );

    \I__5022\ : Span4Mux_h
    port map (
            O => \N__31341\,
            I => \N__31335\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__31338\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_22\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__31335\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_22\
        );

    \I__5019\ : InMux
    port map (
            O => \N__31330\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_21\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__31327\,
            I => \N__31323\
        );

    \I__5017\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31318\
        );

    \I__5016\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31318\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__31318\,
            I => \N__31314\
        );

    \I__5014\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31311\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__31314\,
            I => \N__31308\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__31311\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_23\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__31308\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_23\
        );

    \I__5010\ : InMux
    port map (
            O => \N__31303\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_22\
        );

    \I__5009\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31297\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31293\
        );

    \I__5007\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31290\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__31293\,
            I => \N__31287\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__31290\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_7\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__31287\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_7\
        );

    \I__5003\ : InMux
    port map (
            O => \N__31282\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_6\
        );

    \I__5002\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31276\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31272\
        );

    \I__5000\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31269\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__31272\,
            I => \N__31266\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__31269\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_8\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__31266\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_8\
        );

    \I__4996\ : InMux
    port map (
            O => \N__31261\,
            I => \bfn_11_10_0_\
        );

    \I__4995\ : InMux
    port map (
            O => \N__31258\,
            I => \N__31254\
        );

    \I__4994\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31251\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31248\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__31251\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_9\
        );

    \I__4991\ : Odrv12
    port map (
            O => \N__31248\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_9\
        );

    \I__4990\ : InMux
    port map (
            O => \N__31243\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_8\
        );

    \I__4989\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31236\
        );

    \I__4988\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31233\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31230\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__31233\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_10\
        );

    \I__4985\ : Odrv12
    port map (
            O => \N__31230\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_10\
        );

    \I__4984\ : InMux
    port map (
            O => \N__31225\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_9\
        );

    \I__4983\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31218\
        );

    \I__4982\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31215\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__31218\,
            I => \N__31212\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__31215\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_11\
        );

    \I__4979\ : Odrv12
    port map (
            O => \N__31212\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_11\
        );

    \I__4978\ : InMux
    port map (
            O => \N__31207\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_10\
        );

    \I__4977\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31200\
        );

    \I__4976\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31197\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31194\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__31197\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_12\
        );

    \I__4973\ : Odrv12
    port map (
            O => \N__31194\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_12\
        );

    \I__4972\ : InMux
    port map (
            O => \N__31189\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_11\
        );

    \I__4971\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31183\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31179\
        );

    \I__4969\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31176\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__31179\,
            I => \N__31173\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__31176\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_13\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__31173\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_13\
        );

    \I__4965\ : InMux
    port map (
            O => \N__31168\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_12\
        );

    \I__4964\ : InMux
    port map (
            O => \N__31165\,
            I => \N__31161\
        );

    \I__4963\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31158\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__31161\,
            I => \N__31155\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__31158\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_14\
        );

    \I__4960\ : Odrv12
    port map (
            O => \N__31155\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_14\
        );

    \I__4959\ : InMux
    port map (
            O => \N__31150\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_13\
        );

    \I__4958\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31144\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__31144\,
            I => \N__31140\
        );

    \I__4956\ : InMux
    port map (
            O => \N__31143\,
            I => \N__31137\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__31140\,
            I => \N__31134\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__31137\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_15\
        );

    \I__4953\ : Odrv4
    port map (
            O => \N__31134\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_15\
        );

    \I__4952\ : InMux
    port map (
            O => \N__31129\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_14\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__31126\,
            I => \N__31123\
        );

    \I__4950\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31120\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__31120\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\
        );

    \I__4948\ : CascadeMux
    port map (
            O => \N__31117\,
            I => \N__31113\
        );

    \I__4947\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31110\
        );

    \I__4946\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31107\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__31110\,
            I => \phase_controller_inst2.stoper_hc.counter\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__31107\,
            I => \phase_controller_inst2.stoper_hc.counter\
        );

    \I__4943\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31098\
        );

    \I__4942\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31095\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__31098\,
            I => \N__31092\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__31095\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_0\
        );

    \I__4939\ : Odrv12
    port map (
            O => \N__31092\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_0\
        );

    \I__4938\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31084\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__31084\,
            I => \N__31080\
        );

    \I__4936\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31077\
        );

    \I__4935\ : Span4Mux_v
    port map (
            O => \N__31080\,
            I => \N__31074\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__31077\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_1\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__31074\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_1\
        );

    \I__4932\ : InMux
    port map (
            O => \N__31069\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_0\
        );

    \I__4931\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31062\
        );

    \I__4930\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31059\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31056\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__31059\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_2\
        );

    \I__4927\ : Odrv12
    port map (
            O => \N__31056\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_2\
        );

    \I__4926\ : InMux
    port map (
            O => \N__31051\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_1\
        );

    \I__4925\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31044\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__31047\,
            I => \N__31041\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31038\
        );

    \I__4922\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31035\
        );

    \I__4921\ : Span4Mux_h
    port map (
            O => \N__31038\,
            I => \N__31032\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__31035\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_3\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__31032\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_3\
        );

    \I__4918\ : InMux
    port map (
            O => \N__31027\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_2\
        );

    \I__4917\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31020\
        );

    \I__4916\ : InMux
    port map (
            O => \N__31023\,
            I => \N__31017\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__31020\,
            I => \N__31014\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__31017\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_4\
        );

    \I__4913\ : Odrv12
    port map (
            O => \N__31014\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_4\
        );

    \I__4912\ : InMux
    port map (
            O => \N__31009\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_3\
        );

    \I__4911\ : InMux
    port map (
            O => \N__31006\,
            I => \N__31002\
        );

    \I__4910\ : InMux
    port map (
            O => \N__31005\,
            I => \N__30999\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__31002\,
            I => \N__30996\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__30999\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_5\
        );

    \I__4907\ : Odrv12
    port map (
            O => \N__30996\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_5\
        );

    \I__4906\ : InMux
    port map (
            O => \N__30991\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_4\
        );

    \I__4905\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30984\
        );

    \I__4904\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30981\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30978\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__30981\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_6\
        );

    \I__4901\ : Odrv12
    port map (
            O => \N__30978\,
            I => \phase_controller_inst2.stoper_hc.counterZ0Z_6\
        );

    \I__4900\ : InMux
    port map (
            O => \N__30973\,
            I => \phase_controller_inst2.stoper_hc.counter_cry_5\
        );

    \I__4899\ : InMux
    port map (
            O => \N__30970\,
            I => \bfn_11_8_0_\
        );

    \I__4898\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30964\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__30964\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt20\
        );

    \I__4896\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30958\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__30958\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt18\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__30955\,
            I => \N__30951\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__30954\,
            I => \N__30948\
        );

    \I__4892\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30945\
        );

    \I__4891\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30942\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30939\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30935\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__30939\,
            I => \N__30932\
        );

    \I__4887\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30929\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__30935\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__30932\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__30929\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__30922\,
            I => \N__30919\
        );

    \I__4882\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30916\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__30916\,
            I => \phase_controller_inst2.stoper_hc.un6_running_lt22\
        );

    \I__4880\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30910\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__30910\,
            I => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__4877\ : InMux
    port map (
            O => \N__30904\,
            I => \N__30901\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__30901\,
            I => \phase_controller_inst2.stoper_hc.counter_i_13\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__30898\,
            I => \N__30895\
        );

    \I__4874\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30892\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30889\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__30889\,
            I => \phase_controller_inst2.stoper_hc.counter_i_14\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__30886\,
            I => \N__30883\
        );

    \I__4870\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30880\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__30880\,
            I => \phase_controller_inst2.stoper_hc.counter_i_15\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__30877\,
            I => \N__30874\
        );

    \I__4867\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30871\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__30871\,
            I => \phase_controller_inst2.stoper_hc.counter_i_5\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__30868\,
            I => \N__30865\
        );

    \I__4864\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30862\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__30862\,
            I => \phase_controller_inst2.stoper_hc.counter_i_6\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__4861\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30853\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__30853\,
            I => \phase_controller_inst2.stoper_hc.counter_i_7\
        );

    \I__4859\ : InMux
    port map (
            O => \N__30850\,
            I => \N__30847\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__30847\,
            I => \phase_controller_inst2.stoper_hc.counter_i_8\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__30844\,
            I => \N__30841\
        );

    \I__4856\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30838\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__30838\,
            I => \phase_controller_inst2.stoper_hc.counter_i_9\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__30835\,
            I => \N__30832\
        );

    \I__4853\ : InMux
    port map (
            O => \N__30832\,
            I => \N__30829\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__30829\,
            I => \phase_controller_inst2.stoper_hc.counter_i_10\
        );

    \I__4851\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30823\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__30823\,
            I => \phase_controller_inst2.stoper_hc.counter_i_11\
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__30820\,
            I => \N__30817\
        );

    \I__4848\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30814\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__30814\,
            I => \N__30811\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__30811\,
            I => \phase_controller_inst2.stoper_hc.counter_i_12\
        );

    \I__4845\ : InMux
    port map (
            O => \N__30808\,
            I => \N__30805\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__30805\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__4843\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30799\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__30799\,
            I => \N__30796\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__30796\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__4840\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30790\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__30790\,
            I => \N__30787\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__30787\,
            I => \N__30784\
        );

    \I__4837\ : Sp12to4
    port map (
            O => \N__30784\,
            I => \N__30781\
        );

    \I__4836\ : Span12Mux_s6_v
    port map (
            O => \N__30781\,
            I => \N__30778\
        );

    \I__4835\ : Odrv12
    port map (
            O => \N__30778\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__4834\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30761\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__30774\,
            I => \N__30758\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__30773\,
            I => \N__30755\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__30772\,
            I => \N__30752\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__30771\,
            I => \N__30749\
        );

    \I__4829\ : CascadeMux
    port map (
            O => \N__30770\,
            I => \N__30746\
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__30769\,
            I => \N__30743\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30740\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__30767\,
            I => \N__30737\
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__30766\,
            I => \N__30734\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__30765\,
            I => \N__30731\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__30764\,
            I => \N__30728\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__30761\,
            I => \N__30725\
        );

    \I__4821\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30718\
        );

    \I__4820\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30718\
        );

    \I__4819\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30718\
        );

    \I__4818\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30709\
        );

    \I__4817\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30709\
        );

    \I__4816\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30709\
        );

    \I__4815\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30709\
        );

    \I__4814\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30704\
        );

    \I__4813\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30704\
        );

    \I__4812\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30699\
        );

    \I__4811\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30699\
        );

    \I__4810\ : Span4Mux_v
    port map (
            O => \N__30725\,
            I => \N__30696\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__30718\,
            I => \N__30687\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__30709\,
            I => \N__30687\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30687\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__30699\,
            I => \N__30687\
        );

    \I__4805\ : Span4Mux_v
    port map (
            O => \N__30696\,
            I => \N__30684\
        );

    \I__4804\ : Span4Mux_v
    port map (
            O => \N__30687\,
            I => \N__30681\
        );

    \I__4803\ : Sp12to4
    port map (
            O => \N__30684\,
            I => \N__30676\
        );

    \I__4802\ : Sp12to4
    port map (
            O => \N__30681\,
            I => \N__30676\
        );

    \I__4801\ : Span12Mux_h
    port map (
            O => \N__30676\,
            I => \N__30673\
        );

    \I__4800\ : Odrv12
    port map (
            O => \N__30673\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__30670\,
            I => \N__30667\
        );

    \I__4798\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30664\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30661\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__30661\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__30658\,
            I => \N__30655\
        );

    \I__4794\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30652\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__30652\,
            I => \phase_controller_inst2.stoper_hc.counter_i_0\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__30649\,
            I => \N__30646\
        );

    \I__4791\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30643\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__30643\,
            I => \phase_controller_inst2.stoper_hc.counter_i_1\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__30640\,
            I => \N__30637\
        );

    \I__4788\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30634\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__30634\,
            I => \N__30631\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__30631\,
            I => \phase_controller_inst2.stoper_hc.counter_i_2\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__30628\,
            I => \N__30625\
        );

    \I__4784\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30622\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__30622\,
            I => \phase_controller_inst2.stoper_hc.counter_i_3\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__30619\,
            I => \N__30616\
        );

    \I__4781\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30613\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__30613\,
            I => \N__30610\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__30610\,
            I => \phase_controller_inst2.stoper_hc.counter_i_4\
        );

    \I__4778\ : InMux
    port map (
            O => \N__30607\,
            I => \N__30604\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__30604\,
            I => \N__30601\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__30601\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__4775\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30595\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__30595\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__4773\ : InMux
    port map (
            O => \N__30592\,
            I => \N__30589\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__30589\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__4771\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30583\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__30583\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__4769\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30577\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__30577\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__4767\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30571\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__30571\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__4765\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30565\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__30565\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4763\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30559\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__30559\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__4761\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30553\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__30553\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__4759\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30547\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__30547\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\
        );

    \I__4757\ : InMux
    port map (
            O => \N__30544\,
            I => \N__30541\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__30541\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4755\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30535\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__30535\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__4753\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30529\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__30529\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__4751\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30523\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__30523\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\
        );

    \I__4749\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30517\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__30517\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__4747\ : InMux
    port map (
            O => \N__30514\,
            I => \N__30511\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__30511\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__4745\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30505\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__30505\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__4743\ : InMux
    port map (
            O => \N__30502\,
            I => \bfn_10_17_0_\
        );

    \I__4742\ : IoInMux
    port map (
            O => \N__30499\,
            I => \N__30496\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30493\
        );

    \I__4740\ : Span4Mux_s2_v
    port map (
            O => \N__30493\,
            I => \N__30490\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__30490\,
            I => \N__30487\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__30487\,
            I => \N__30484\
        );

    \I__4737\ : Span4Mux_v
    port map (
            O => \N__30484\,
            I => \N__30481\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__30481\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__4735\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30475\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__30475\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__4733\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30469\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__30469\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__30466\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__4730\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30460\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__30460\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__30457\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_cascade_\
        );

    \I__4727\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30451\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__30451\,
            I => \N__30448\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__30448\,
            I => \N__30445\
        );

    \I__4724\ : Span4Mux_h
    port map (
            O => \N__30445\,
            I => \N__30442\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__30442\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__30439\,
            I => \N__30436\
        );

    \I__4721\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30433\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30430\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__30430\,
            I => \N__30427\
        );

    \I__4718\ : Span4Mux_h
    port map (
            O => \N__30427\,
            I => \N__30424\
        );

    \I__4717\ : Odrv4
    port map (
            O => \N__30424\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt16\
        );

    \I__4716\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30418\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30415\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__30415\,
            I => \N__30412\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__30412\,
            I => \N__30409\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__30409\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\
        );

    \I__4711\ : CascadeMux
    port map (
            O => \N__30406\,
            I => \N__30403\
        );

    \I__4710\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30400\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__30400\,
            I => \N__30397\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__30397\,
            I => \N__30394\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__30394\,
            I => \N__30391\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__30391\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt18\
        );

    \I__4705\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30385\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__30385\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__30382\,
            I => \N__30379\
        );

    \I__4702\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30376\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__30376\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt24\
        );

    \I__4700\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30370\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__30370\,
            I => \phase_controller_inst1.stoper_tr.un6_running_lt26\
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__30367\,
            I => \N__30364\
        );

    \I__4697\ : InMux
    port map (
            O => \N__30364\,
            I => \N__30361\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__30361\,
            I => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\
        );

    \I__4695\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30355\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__30355\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__30352\,
            I => \N__30349\
        );

    \I__4692\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30346\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30343\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__30343\,
            I => \phase_controller_inst1.stoper_tr.counter_i_7\
        );

    \I__4689\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30337\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__30337\,
            I => \phase_controller_inst1.stoper_tr.counter_i_8\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__4686\ : InMux
    port map (
            O => \N__30331\,
            I => \N__30328\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__30328\,
            I => \phase_controller_inst1.stoper_tr.counter_i_9\
        );

    \I__4684\ : InMux
    port map (
            O => \N__30325\,
            I => \N__30322\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__30322\,
            I => \phase_controller_inst1.stoper_tr.counter_i_10\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__30319\,
            I => \N__30316\
        );

    \I__4681\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30313\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__30313\,
            I => \phase_controller_inst1.stoper_tr.counter_i_11\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__30310\,
            I => \N__30307\
        );

    \I__4678\ : InMux
    port map (
            O => \N__30307\,
            I => \N__30304\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__30304\,
            I => \phase_controller_inst1.stoper_tr.counter_i_12\
        );

    \I__4676\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30298\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__30298\,
            I => \N__30295\
        );

    \I__4674\ : Odrv12
    port map (
            O => \N__30295\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__30292\,
            I => \N__30289\
        );

    \I__4672\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30286\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__30286\,
            I => \phase_controller_inst1.stoper_tr.counter_i_13\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__30283\,
            I => \N__30280\
        );

    \I__4669\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30277\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__30277\,
            I => \phase_controller_inst1.stoper_tr.counter_i_14\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30271\
        );

    \I__4666\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30268\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__30268\,
            I => \phase_controller_inst1.stoper_tr.counter_i_15\
        );

    \I__4664\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30261\
        );

    \I__4663\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30258\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30255\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__30258\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_3
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__30255\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_3
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__30250\,
            I => \N__30247\
        );

    \I__4658\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30244\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__30244\,
            I => \phase_controller_inst1.stoper_tr.counter_i_0\
        );

    \I__4656\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30238\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__30238\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__30235\,
            I => \N__30232\
        );

    \I__4653\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30229\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__30229\,
            I => \phase_controller_inst1.stoper_tr.counter_i_1\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__4650\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__30220\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\
        );

    \I__4648\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30214\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__30214\,
            I => \phase_controller_inst1.stoper_tr.counter_i_2\
        );

    \I__4646\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30208\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__30208\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__4643\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30199\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__30199\,
            I => \phase_controller_inst1.stoper_tr.counter_i_3\
        );

    \I__4641\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__30193\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__30190\,
            I => \N__30187\
        );

    \I__4638\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30184\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__30184\,
            I => \phase_controller_inst1.stoper_tr.counter_i_4\
        );

    \I__4636\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__30178\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__30175\,
            I => \N__30172\
        );

    \I__4633\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30169\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__30169\,
            I => \phase_controller_inst1.stoper_tr.counter_i_5\
        );

    \I__4631\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30163\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__30163\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__30160\,
            I => \N__30157\
        );

    \I__4628\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__30154\,
            I => \phase_controller_inst1.stoper_tr.counter_i_6\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__30151\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\
        );

    \I__4625\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30145\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__30145\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\
        );

    \I__4623\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30138\
        );

    \I__4622\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30135\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__30138\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__30135\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__4619\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30127\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30124\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__30124\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\
        );

    \I__4616\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30117\
        );

    \I__4615\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30114\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__30117\,
            I => \N__30111\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__30114\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_1
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__30111\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_1
        );

    \I__4611\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30102\
        );

    \I__4610\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30099\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30096\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__30099\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_6
        );

    \I__4607\ : Odrv4
    port map (
            O => \N__30096\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_6
        );

    \I__4606\ : InMux
    port map (
            O => \N__30091\,
            I => \N__30087\
        );

    \I__4605\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30084\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__30087\,
            I => \N__30081\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__30084\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_5
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__30081\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_5
        );

    \I__4601\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30073\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__30073\,
            I => \N__30070\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__30070\,
            I => \N__30066\
        );

    \I__4598\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30063\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__30066\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_13
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__30063\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_13
        );

    \I__4595\ : InMux
    port map (
            O => \N__30058\,
            I => \N__30054\
        );

    \I__4594\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30051\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__30054\,
            I => \N__30048\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__30051\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_7
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__30048\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_7
        );

    \I__4590\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30039\
        );

    \I__4589\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30036\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__30039\,
            I => \N__30033\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__30036\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_4
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__30033\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_4
        );

    \I__4585\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30025\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__30025\,
            I => \N__30021\
        );

    \I__4583\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30018\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__30021\,
            I => \N__30013\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__30018\,
            I => \N__30013\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__30013\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_2
        );

    \I__4579\ : InMux
    port map (
            O => \N__30010\,
            I => \N__30007\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__30007\,
            I => \N__30004\
        );

    \I__4577\ : Span4Mux_v
    port map (
            O => \N__30004\,
            I => \N__30000\
        );

    \I__4576\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29997\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__30000\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__29997\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4573\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29985\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__29988\,
            I => \N__29982\
        );

    \I__4570\ : Span4Mux_h
    port map (
            O => \N__29985\,
            I => \N__29979\
        );

    \I__4569\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29976\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__29979\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__29976\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4566\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29967\
        );

    \I__4565\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29964\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__29967\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__29964\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4562\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29956\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__29956\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\
        );

    \I__4560\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29949\
        );

    \I__4559\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29946\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__29949\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__29946\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4556\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29938\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__29938\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\
        );

    \I__4554\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29931\
        );

    \I__4553\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29928\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29923\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__29928\,
            I => \N__29923\
        );

    \I__4550\ : Span4Mux_v
    port map (
            O => \N__29923\,
            I => \N__29920\
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__29920\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__4548\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29914\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__29914\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__29911\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\
        );

    \I__4545\ : InMux
    port map (
            O => \N__29908\,
            I => \N__29905\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__29905\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\
        );

    \I__4543\ : InMux
    port map (
            O => \N__29902\,
            I => \N__29898\
        );

    \I__4542\ : InMux
    port map (
            O => \N__29901\,
            I => \N__29895\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__29898\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__29895\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__4539\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29887\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__29887\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\
        );

    \I__4537\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29881\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29877\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__29880\,
            I => \N__29874\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__29877\,
            I => \N__29871\
        );

    \I__4533\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29868\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__29871\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__29868\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__4530\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29860\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__29860\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__4528\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29854\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__29854\,
            I => \N__29851\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__29851\,
            I => \N__29847\
        );

    \I__4525\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29844\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__29847\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__29844\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__4522\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29836\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__29836\,
            I => \N__29832\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__29835\,
            I => \N__29829\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__29832\,
            I => \N__29825\
        );

    \I__4518\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29822\
        );

    \I__4517\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29819\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__29825\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__29822\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__29819\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__29812\,
            I => \N__29809\
        );

    \I__4512\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29805\
        );

    \I__4511\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29802\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__29805\,
            I => \N__29799\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__29802\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4508\ : Odrv4
    port map (
            O => \N__29799\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__4507\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29791\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__29791\,
            I => \N__29787\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__29790\,
            I => \N__29784\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29780\
        );

    \I__4503\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29777\
        );

    \I__4502\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29774\
        );

    \I__4501\ : Odrv4
    port map (
            O => \N__29780\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__29777\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__29774\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__4498\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29763\
        );

    \I__4497\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29760\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__29763\,
            I => \N__29757\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__29760\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__29757\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4493\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29748\
        );

    \I__4492\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29745\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__29748\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__29745\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4489\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29736\
        );

    \I__4488\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29733\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__29736\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__29733\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__4485\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29725\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__29725\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\
        );

    \I__4483\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29719\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N__29716\
        );

    \I__4481\ : Span4Mux_h
    port map (
            O => \N__29716\,
            I => \N__29712\
        );

    \I__4480\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29709\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__29712\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__29709\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4477\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29701\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29698\
        );

    \I__4475\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29694\
        );

    \I__4474\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29691\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__29694\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__29691\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4471\ : InMux
    port map (
            O => \N__29686\,
            I => \N__29683\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__29683\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\
        );

    \I__4468\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29674\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__29674\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\
        );

    \I__4466\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29668\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29665\
        );

    \I__4464\ : Span4Mux_h
    port map (
            O => \N__29665\,
            I => \N__29661\
        );

    \I__4463\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29658\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__29661\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__29658\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4460\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29648\
        );

    \I__4459\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29643\
        );

    \I__4458\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29643\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__29648\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__29643\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__4455\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29635\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__29635\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__29632\,
            I => \N__29629\
        );

    \I__4452\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29625\
        );

    \I__4451\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29622\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29619\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29616\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__29619\,
            I => \N__29613\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__29616\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__29613\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__4445\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29605\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__29605\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__4443\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29599\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__29599\,
            I => \N__29595\
        );

    \I__4441\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29592\
        );

    \I__4440\ : Span4Mux_h
    port map (
            O => \N__29595\,
            I => \N__29589\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__29592\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__29589\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4437\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29581\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__29581\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__29578\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__4434\ : InMux
    port map (
            O => \N__29575\,
            I => \N__29572\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__29572\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__29569\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__4431\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29562\
        );

    \I__4430\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29559\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__29562\,
            I => \N__29556\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__29559\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__29556\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__4426\ : InMux
    port map (
            O => \N__29551\,
            I => \N__29548\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__29548\,
            I => \N__29545\
        );

    \I__4424\ : Span4Mux_v
    port map (
            O => \N__29545\,
            I => \N__29542\
        );

    \I__4423\ : Odrv4
    port map (
            O => \N__29542\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\
        );

    \I__4422\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29536\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__29536\,
            I => \N__29532\
        );

    \I__4420\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29529\
        );

    \I__4419\ : Odrv4
    port map (
            O => \N__29532\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__29529\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__4417\ : InMux
    port map (
            O => \N__29524\,
            I => \N__29518\
        );

    \I__4416\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29518\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__29518\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__4414\ : InMux
    port map (
            O => \N__29515\,
            I => \N__29512\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__29512\,
            I => \N__29508\
        );

    \I__4412\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29505\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__29508\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__29505\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__4409\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29497\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__29497\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__29494\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\
        );

    \I__4406\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29488\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__29488\,
            I => \N__29485\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__29485\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\
        );

    \I__4403\ : IoInMux
    port map (
            O => \N__29482\,
            I => \N__29479\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__29479\,
            I => \N__29476\
        );

    \I__4401\ : Span4Mux_s0_v
    port map (
            O => \N__29476\,
            I => \N__29473\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__29473\,
            I => \N__29470\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__29470\,
            I => s4_phy_c
        );

    \I__4398\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29462\
        );

    \I__4397\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29459\
        );

    \I__4396\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29456\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29451\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29451\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__29456\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__29451\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4391\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29443\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__29443\,
            I => \N__29438\
        );

    \I__4389\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29433\
        );

    \I__4388\ : InMux
    port map (
            O => \N__29441\,
            I => \N__29433\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__29438\,
            I => \N__29428\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__29433\,
            I => \N__29428\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__29428\,
            I => \N__29425\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__29425\,
            I => \N__29422\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__29422\,
            I => il_min_comp2_c
        );

    \I__4382\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29416\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__29416\,
            I => \N__29413\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__29413\,
            I => \N__29410\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__29410\,
            I => \N__29406\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__29409\,
            I => \N__29401\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__29406\,
            I => \N__29398\
        );

    \I__4376\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29395\
        );

    \I__4375\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29390\
        );

    \I__4374\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29390\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__29398\,
            I => \N__29387\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__29395\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__29390\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__29387\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__4369\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29377\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__29377\,
            I => \N__29372\
        );

    \I__4367\ : InMux
    port map (
            O => \N__29376\,
            I => \N__29367\
        );

    \I__4366\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29367\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__29372\,
            I => \N__29362\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__29367\,
            I => \N__29362\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__29362\,
            I => \N__29359\
        );

    \I__4362\ : IoSpan4Mux
    port map (
            O => \N__29359\,
            I => \N__29356\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__29356\,
            I => il_max_comp2_c
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__29353\,
            I => \N__29350\
        );

    \I__4359\ : InMux
    port map (
            O => \N__29350\,
            I => \N__29346\
        );

    \I__4358\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29343\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__29346\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__29343\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__29338\,
            I => \phase_controller_inst2.state_ns_0_0_1_cascade_\
        );

    \I__4354\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29332\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__29332\,
            I => \N__29328\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__29331\,
            I => \N__29324\
        );

    \I__4351\ : Sp12to4
    port map (
            O => \N__29328\,
            I => \N__29320\
        );

    \I__4350\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29315\
        );

    \I__4349\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29315\
        );

    \I__4348\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29312\
        );

    \I__4347\ : Span12Mux_v
    port map (
            O => \N__29320\,
            I => \N__29309\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__29315\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__29312\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4344\ : Odrv12
    port map (
            O => \N__29309\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__29302\,
            I => \phase_controller_inst2.stoper_tr.un4_start_0_cascade_\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__29299\,
            I => \N__29294\
        );

    \I__4341\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29291\
        );

    \I__4340\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29286\
        );

    \I__4339\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29286\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__29291\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__29286\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__4336\ : IoInMux
    port map (
            O => \N__29281\,
            I => \N__29278\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__29278\,
            I => \N__29275\
        );

    \I__4334\ : Span12Mux_s6_v
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__4333\ : Odrv12
    port map (
            O => \N__29272\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__4332\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29261\
        );

    \I__4331\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29258\
        );

    \I__4330\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29255\
        );

    \I__4329\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29248\
        );

    \I__4328\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29248\
        );

    \I__4327\ : InMux
    port map (
            O => \N__29264\,
            I => \N__29248\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__29261\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__29258\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__29255\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__29248\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__4322\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29233\
        );

    \I__4321\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29233\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29230\
        );

    \I__4319\ : Span4Mux_v
    port map (
            O => \N__29230\,
            I => \N__29227\
        );

    \I__4318\ : Span4Mux_v
    port map (
            O => \N__29227\,
            I => \N__29224\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__29224\,
            I => \N__29221\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__29221\,
            I => \N__29217\
        );

    \I__4315\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29214\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__29217\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__29214\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__29209\,
            I => \N__29206\
        );

    \I__4311\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29203\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__29203\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__4309\ : InMux
    port map (
            O => \N__29200\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__4308\ : InMux
    port map (
            O => \N__29197\,
            I => \N__29194\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__29194\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__4306\ : InMux
    port map (
            O => \N__29191\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__4305\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29185\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__29185\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__4303\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29179\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__29179\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__4301\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29173\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__29173\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4299\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29167\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__29167\,
            I => \N__29164\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__29164\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__4296\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29158\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__29158\,
            I => \N__29155\
        );

    \I__4294\ : Odrv12
    port map (
            O => \N__29155\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__4293\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29149\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__29149\,
            I => \N__29146\
        );

    \I__4291\ : Odrv12
    port map (
            O => \N__29146\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__4290\ : IoInMux
    port map (
            O => \N__29143\,
            I => \N__29140\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__29140\,
            I => \N__29137\
        );

    \I__4288\ : Span4Mux_s3_v
    port map (
            O => \N__29137\,
            I => \N__29134\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__29134\,
            I => s3_phy_c
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__29131\,
            I => \N__29128\
        );

    \I__4285\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29125\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__29125\,
            I => \N__29122\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__29122\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__4282\ : InMux
    port map (
            O => \N__29119\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__4281\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29113\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__29113\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__4279\ : InMux
    port map (
            O => \N__29110\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__29107\,
            I => \N__29104\
        );

    \I__4277\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29101\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__29101\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__4275\ : InMux
    port map (
            O => \N__29098\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__29095\,
            I => \N__29092\
        );

    \I__4273\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29089\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29086\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__29083\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__4269\ : InMux
    port map (
            O => \N__29080\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__29077\,
            I => \N__29074\
        );

    \I__4267\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29071\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__29071\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__4265\ : InMux
    port map (
            O => \N__29068\,
            I => \bfn_9_21_0_\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__4263\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29059\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__29059\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__4261\ : InMux
    port map (
            O => \N__29056\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__4260\ : CascadeMux
    port map (
            O => \N__29053\,
            I => \N__29050\
        );

    \I__4259\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29047\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__29047\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__4257\ : InMux
    port map (
            O => \N__29044\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__29041\,
            I => \N__29038\
        );

    \I__4255\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29035\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__29035\,
            I => \N__29032\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__29032\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__4252\ : InMux
    port map (
            O => \N__29029\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__29026\,
            I => \N__29023\
        );

    \I__4250\ : InMux
    port map (
            O => \N__29023\,
            I => \N__29020\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__29020\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__4248\ : InMux
    port map (
            O => \N__29017\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__29014\,
            I => \N__29011\
        );

    \I__4246\ : InMux
    port map (
            O => \N__29011\,
            I => \N__29008\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__29008\,
            I => \N__29005\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__4243\ : Sp12to4
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__4242\ : Span12Mux_h
    port map (
            O => \N__28999\,
            I => \N__28996\
        );

    \I__4241\ : Span12Mux_v
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__4240\ : Odrv12
    port map (
            O => \N__28993\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__4239\ : InMux
    port map (
            O => \N__28990\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__4237\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28981\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__28981\,
            I => \N__28978\
        );

    \I__4235\ : Span4Mux_h
    port map (
            O => \N__28978\,
            I => \N__28975\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__4233\ : Sp12to4
    port map (
            O => \N__28972\,
            I => \N__28969\
        );

    \I__4232\ : Span12Mux_v
    port map (
            O => \N__28969\,
            I => \N__28966\
        );

    \I__4231\ : Odrv12
    port map (
            O => \N__28966\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__4230\ : InMux
    port map (
            O => \N__28963\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__28960\,
            I => \N__28957\
        );

    \I__4228\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28954\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28951\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__28951\,
            I => \N__28948\
        );

    \I__4225\ : Sp12to4
    port map (
            O => \N__28948\,
            I => \N__28945\
        );

    \I__4224\ : Span12Mux_v
    port map (
            O => \N__28945\,
            I => \N__28942\
        );

    \I__4223\ : Odrv12
    port map (
            O => \N__28942\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__4222\ : InMux
    port map (
            O => \N__28939\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__28936\,
            I => \N__28933\
        );

    \I__4220\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28930\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__28930\,
            I => \N__28927\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__28927\,
            I => \N__28924\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__28924\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__4216\ : InMux
    port map (
            O => \N__28921\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__4215\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28915\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__28915\,
            I => \N__28912\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__28912\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__4212\ : InMux
    port map (
            O => \N__28909\,
            I => \bfn_9_20_0_\
        );

    \I__4211\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28903\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__28903\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__4209\ : InMux
    port map (
            O => \N__28900\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__28897\,
            I => \N__28894\
        );

    \I__4207\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28891\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__28891\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__4205\ : InMux
    port map (
            O => \N__28888\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__4204\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28882\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__28882\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__4202\ : InMux
    port map (
            O => \N__28879\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__4200\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28870\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28867\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__28867\,
            I => \N__28864\
        );

    \I__4197\ : Sp12to4
    port map (
            O => \N__28864\,
            I => \N__28861\
        );

    \I__4196\ : Span12Mux_h
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__4195\ : Span12Mux_v
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__4194\ : Odrv12
    port map (
            O => \N__28855\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__4193\ : InMux
    port map (
            O => \N__28852\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__4191\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28843\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__28843\,
            I => \N__28840\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__28840\,
            I => \N__28837\
        );

    \I__4188\ : Sp12to4
    port map (
            O => \N__28837\,
            I => \N__28834\
        );

    \I__4187\ : Span12Mux_v
    port map (
            O => \N__28834\,
            I => \N__28831\
        );

    \I__4186\ : Odrv12
    port map (
            O => \N__28831\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__4185\ : InMux
    port map (
            O => \N__28828\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__28825\,
            I => \N__28822\
        );

    \I__4183\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28816\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__28816\,
            I => \N__28813\
        );

    \I__4180\ : Sp12to4
    port map (
            O => \N__28813\,
            I => \N__28810\
        );

    \I__4179\ : Span12Mux_v
    port map (
            O => \N__28810\,
            I => \N__28807\
        );

    \I__4178\ : Odrv12
    port map (
            O => \N__28807\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__4177\ : InMux
    port map (
            O => \N__28804\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__28801\,
            I => \N__28798\
        );

    \I__4175\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28795\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28792\
        );

    \I__4173\ : Sp12to4
    port map (
            O => \N__28792\,
            I => \N__28789\
        );

    \I__4172\ : Span12Mux_v
    port map (
            O => \N__28789\,
            I => \N__28786\
        );

    \I__4171\ : Odrv12
    port map (
            O => \N__28786\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__4170\ : InMux
    port map (
            O => \N__28783\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__4169\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28777\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28774\
        );

    \I__4167\ : Span4Mux_v
    port map (
            O => \N__28774\,
            I => \N__28771\
        );

    \I__4166\ : Sp12to4
    port map (
            O => \N__28771\,
            I => \N__28768\
        );

    \I__4165\ : Span12Mux_h
    port map (
            O => \N__28768\,
            I => \N__28765\
        );

    \I__4164\ : Span12Mux_v
    port map (
            O => \N__28765\,
            I => \N__28762\
        );

    \I__4163\ : Odrv12
    port map (
            O => \N__28762\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__4162\ : InMux
    port map (
            O => \N__28759\,
            I => \bfn_9_19_0_\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__28756\,
            I => \N__28753\
        );

    \I__4160\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__4158\ : Span12Mux_h
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__4157\ : Span12Mux_v
    port map (
            O => \N__28744\,
            I => \N__28741\
        );

    \I__4156\ : Odrv12
    port map (
            O => \N__28741\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__4155\ : InMux
    port map (
            O => \N__28738\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__28735\,
            I => \N__28732\
        );

    \I__4153\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28729\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__28729\,
            I => \N__28726\
        );

    \I__4151\ : Span4Mux_v
    port map (
            O => \N__28726\,
            I => \N__28723\
        );

    \I__4150\ : Sp12to4
    port map (
            O => \N__28723\,
            I => \N__28720\
        );

    \I__4149\ : Span12Mux_h
    port map (
            O => \N__28720\,
            I => \N__28717\
        );

    \I__4148\ : Odrv12
    port map (
            O => \N__28717\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__4147\ : InMux
    port map (
            O => \N__28714\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__28711\,
            I => \N__28708\
        );

    \I__4145\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28705\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28702\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__28702\,
            I => \N__28699\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__28699\,
            I => \N__28696\
        );

    \I__4141\ : Sp12to4
    port map (
            O => \N__28696\,
            I => \N__28693\
        );

    \I__4140\ : Span12Mux_v
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__28690\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__4138\ : InMux
    port map (
            O => \N__28687\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__4137\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__28681\,
            I => \N__28677\
        );

    \I__4135\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28674\
        );

    \I__4134\ : Odrv12
    port map (
            O => \N__28677\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_25
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__28674\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_25
        );

    \I__4132\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28663\
        );

    \I__4131\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28663\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__28663\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\
        );

    \I__4129\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28657\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__28657\,
            I => \N__28653\
        );

    \I__4127\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28650\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__28653\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_26
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__28650\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_26
        );

    \I__4124\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28639\
        );

    \I__4123\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28639\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__28639\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\
        );

    \I__4121\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28633\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28629\
        );

    \I__4119\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28626\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__28629\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_27
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__28626\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_27
        );

    \I__4116\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28615\
        );

    \I__4115\ : InMux
    port map (
            O => \N__28620\,
            I => \N__28615\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__28615\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__28612\,
            I => \N__28609\
        );

    \I__4112\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28606\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__28606\,
            I => \N__28603\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__4109\ : Sp12to4
    port map (
            O => \N__28600\,
            I => \N__28597\
        );

    \I__4108\ : Span12Mux_h
    port map (
            O => \N__28597\,
            I => \N__28594\
        );

    \I__4107\ : Span12Mux_v
    port map (
            O => \N__28594\,
            I => \N__28591\
        );

    \I__4106\ : Odrv12
    port map (
            O => \N__28591\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__28588\,
            I => \N__28585\
        );

    \I__4104\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__28582\,
            I => \N__28579\
        );

    \I__4102\ : Span4Mux_v
    port map (
            O => \N__28579\,
            I => \N__28576\
        );

    \I__4101\ : Sp12to4
    port map (
            O => \N__28576\,
            I => \N__28573\
        );

    \I__4100\ : Span12Mux_h
    port map (
            O => \N__28573\,
            I => \N__28570\
        );

    \I__4099\ : Odrv12
    port map (
            O => \N__28570\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__4098\ : InMux
    port map (
            O => \N__28567\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__28564\,
            I => \N__28561\
        );

    \I__4096\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28558\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__28558\,
            I => \N__28555\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__28555\,
            I => \N__28552\
        );

    \I__4093\ : Sp12to4
    port map (
            O => \N__28552\,
            I => \N__28549\
        );

    \I__4092\ : Span12Mux_h
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__4091\ : Odrv12
    port map (
            O => \N__28546\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__4090\ : InMux
    port map (
            O => \N__28543\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__4088\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28534\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28531\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__28531\,
            I => \N__28528\
        );

    \I__4085\ : Sp12to4
    port map (
            O => \N__28528\,
            I => \N__28525\
        );

    \I__4084\ : Span12Mux_h
    port map (
            O => \N__28525\,
            I => \N__28522\
        );

    \I__4083\ : Odrv12
    port map (
            O => \N__28522\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__4082\ : InMux
    port map (
            O => \N__28519\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__4081\ : InMux
    port map (
            O => \N__28516\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__4080\ : InMux
    port map (
            O => \N__28513\,
            I => \N__28510\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__28510\,
            I => \N__28507\
        );

    \I__4078\ : Span12Mux_h
    port map (
            O => \N__28507\,
            I => \N__28504\
        );

    \I__4077\ : Odrv12
    port map (
            O => \N__28504\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__4076\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28498\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__28498\,
            I => \N__28495\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__28495\,
            I => \N__28492\
        );

    \I__4073\ : Sp12to4
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__4072\ : Span12Mux_s9_h
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__4071\ : Odrv12
    port map (
            O => \N__28486\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\
        );

    \I__4070\ : InMux
    port map (
            O => \N__28483\,
            I => \bfn_9_16_0_\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__4068\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__28468\,
            I => \N__28465\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__28465\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__4063\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28459\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28456\
        );

    \I__4061\ : Span12Mux_s9_h
    port map (
            O => \N__28456\,
            I => \N__28453\
        );

    \I__4060\ : Odrv12
    port map (
            O => \N__28453\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\
        );

    \I__4059\ : InMux
    port map (
            O => \N__28450\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__4058\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28444\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__28444\,
            I => \N__28441\
        );

    \I__4056\ : Span12Mux_h
    port map (
            O => \N__28441\,
            I => \N__28438\
        );

    \I__4055\ : Odrv12
    port map (
            O => \N__28438\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__4054\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28432\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__28432\,
            I => \N__28429\
        );

    \I__4052\ : Span4Mux_v
    port map (
            O => \N__28429\,
            I => \N__28426\
        );

    \I__4051\ : Sp12to4
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__4050\ : Span12Mux_s9_h
    port map (
            O => \N__28423\,
            I => \N__28420\
        );

    \I__4049\ : Odrv12
    port map (
            O => \N__28420\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\
        );

    \I__4048\ : InMux
    port map (
            O => \N__28417\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__28414\,
            I => \N__28406\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__28413\,
            I => \N__28402\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__28412\,
            I => \N__28398\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__28411\,
            I => \N__28395\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__28410\,
            I => \N__28392\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__28409\,
            I => \N__28389\
        );

    \I__4041\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28385\
        );

    \I__4040\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28376\
        );

    \I__4039\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28376\
        );

    \I__4038\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28376\
        );

    \I__4037\ : InMux
    port map (
            O => \N__28398\,
            I => \N__28376\
        );

    \I__4036\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28373\
        );

    \I__4035\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28366\
        );

    \I__4034\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28366\
        );

    \I__4033\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28366\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28363\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__28376\,
            I => \N__28360\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28355\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__28366\,
            I => \N__28355\
        );

    \I__4028\ : Span12Mux_s10_v
    port map (
            O => \N__28363\,
            I => \N__28352\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__28360\,
            I => \N__28347\
        );

    \I__4026\ : Span4Mux_v
    port map (
            O => \N__28355\,
            I => \N__28347\
        );

    \I__4025\ : Span12Mux_h
    port map (
            O => \N__28352\,
            I => \N__28344\
        );

    \I__4024\ : Sp12to4
    port map (
            O => \N__28347\,
            I => \N__28341\
        );

    \I__4023\ : Span12Mux_h
    port map (
            O => \N__28344\,
            I => \N__28338\
        );

    \I__4022\ : Span12Mux_h
    port map (
            O => \N__28341\,
            I => \N__28335\
        );

    \I__4021\ : Odrv12
    port map (
            O => \N__28338\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__4020\ : Odrv12
    port map (
            O => \N__28335\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__28330\,
            I => \N__28327\
        );

    \I__4018\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28324\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__28324\,
            I => \N__28321\
        );

    \I__4016\ : Span4Mux_h
    port map (
            O => \N__28321\,
            I => \N__28318\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__28318\,
            I => \N__28315\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__28315\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__4013\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28309\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__28309\,
            I => \N__28306\
        );

    \I__4011\ : Sp12to4
    port map (
            O => \N__28306\,
            I => \N__28303\
        );

    \I__4010\ : Span12Mux_v
    port map (
            O => \N__28303\,
            I => \N__28300\
        );

    \I__4009\ : Odrv12
    port map (
            O => \N__28300\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\
        );

    \I__4008\ : InMux
    port map (
            O => \N__28297\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__4007\ : InMux
    port map (
            O => \N__28294\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__4006\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28288\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28285\
        );

    \I__4004\ : Span12Mux_v
    port map (
            O => \N__28285\,
            I => \N__28282\
        );

    \I__4003\ : Odrv12
    port map (
            O => \N__28282\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO\
        );

    \I__4002\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28276\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__28276\,
            I => \N__28272\
        );

    \I__4000\ : InMux
    port map (
            O => \N__28275\,
            I => \N__28269\
        );

    \I__3999\ : Odrv12
    port map (
            O => \N__28272\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_24
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__28269\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_24
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__28264\,
            I => \N__28260\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__28263\,
            I => \N__28257\
        );

    \I__3995\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28252\
        );

    \I__3994\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28252\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__28252\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\
        );

    \I__3992\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28246\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N__28243\
        );

    \I__3990\ : Span12Mux_h
    port map (
            O => \N__28243\,
            I => \N__28240\
        );

    \I__3989\ : Odrv12
    port map (
            O => \N__28240\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__3987\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28231\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__3985\ : Span4Mux_v
    port map (
            O => \N__28228\,
            I => \N__28225\
        );

    \I__3984\ : Span4Mux_h
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__3983\ : Sp12to4
    port map (
            O => \N__28222\,
            I => \N__28219\
        );

    \I__3982\ : Odrv12
    port map (
            O => \N__28219\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__3981\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__28204\,
            I => \N__28201\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__28201\,
            I => \N__28198\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__28198\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_8\
        );

    \I__3974\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28192\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28189\
        );

    \I__3972\ : Span4Mux_h
    port map (
            O => \N__28189\,
            I => \N__28186\
        );

    \I__3971\ : Span4Mux_h
    port map (
            O => \N__28186\,
            I => \N__28183\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__28183\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__28180\,
            I => \N__28177\
        );

    \I__3968\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28174\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__28174\,
            I => \N__28171\
        );

    \I__3966\ : Span4Mux_h
    port map (
            O => \N__28171\,
            I => \N__28168\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__28168\,
            I => \N__28165\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__28165\,
            I => \N__28162\
        );

    \I__3963\ : Span4Mux_h
    port map (
            O => \N__28162\,
            I => \N__28159\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__28159\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__3961\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__28153\,
            I => \N__28150\
        );

    \I__3959\ : Span12Mux_s9_h
    port map (
            O => \N__28150\,
            I => \N__28147\
        );

    \I__3958\ : Odrv12
    port map (
            O => \N__28147\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\
        );

    \I__3957\ : InMux
    port map (
            O => \N__28144\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__3956\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28138\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__3954\ : Span4Mux_v
    port map (
            O => \N__28135\,
            I => \N__28132\
        );

    \I__3953\ : Sp12to4
    port map (
            O => \N__28132\,
            I => \N__28129\
        );

    \I__3952\ : Span12Mux_h
    port map (
            O => \N__28129\,
            I => \N__28126\
        );

    \I__3951\ : Odrv12
    port map (
            O => \N__28126\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__28123\,
            I => \N__28120\
        );

    \I__3949\ : InMux
    port map (
            O => \N__28120\,
            I => \N__28117\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__28117\,
            I => \N__28114\
        );

    \I__3947\ : Span12Mux_h
    port map (
            O => \N__28114\,
            I => \N__28111\
        );

    \I__3946\ : Odrv12
    port map (
            O => \N__28111\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__3945\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28105\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__28105\,
            I => \N__28102\
        );

    \I__3943\ : Span4Mux_v
    port map (
            O => \N__28102\,
            I => \N__28099\
        );

    \I__3942\ : Span4Mux_h
    port map (
            O => \N__28099\,
            I => \N__28096\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__28096\,
            I => \N__28093\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__28090\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\
        );

    \I__3938\ : InMux
    port map (
            O => \N__28087\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__3937\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28081\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__28081\,
            I => \N__28078\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__28078\,
            I => \N__28075\
        );

    \I__3934\ : Sp12to4
    port map (
            O => \N__28075\,
            I => \N__28072\
        );

    \I__3933\ : Span12Mux_h
    port map (
            O => \N__28072\,
            I => \N__28069\
        );

    \I__3932\ : Odrv12
    port map (
            O => \N__28069\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__28066\,
            I => \N__28063\
        );

    \I__3930\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28060\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28057\
        );

    \I__3928\ : Span12Mux_h
    port map (
            O => \N__28057\,
            I => \N__28054\
        );

    \I__3927\ : Odrv12
    port map (
            O => \N__28054\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__3926\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28048\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__28048\,
            I => \N__28045\
        );

    \I__3924\ : Sp12to4
    port map (
            O => \N__28045\,
            I => \N__28042\
        );

    \I__3923\ : Span12Mux_v
    port map (
            O => \N__28042\,
            I => \N__28039\
        );

    \I__3922\ : Odrv12
    port map (
            O => \N__28039\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\
        );

    \I__3921\ : InMux
    port map (
            O => \N__28036\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__28033\,
            I => \N__28030\
        );

    \I__3919\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28027\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__28027\,
            I => \N__28024\
        );

    \I__3917\ : Span4Mux_h
    port map (
            O => \N__28024\,
            I => \N__28021\
        );

    \I__3916\ : Span4Mux_h
    port map (
            O => \N__28021\,
            I => \N__28018\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__28018\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__3914\ : InMux
    port map (
            O => \N__28015\,
            I => \N__28012\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__28012\,
            I => \N__28009\
        );

    \I__3912\ : Span12Mux_v
    port map (
            O => \N__28009\,
            I => \N__28006\
        );

    \I__3911\ : Odrv12
    port map (
            O => \N__28006\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\
        );

    \I__3910\ : InMux
    port map (
            O => \N__28003\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__3909\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27997\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__3907\ : Odrv12
    port map (
            O => \N__27994\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__3906\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27988\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27985\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__27985\,
            I => \N__27982\
        );

    \I__3903\ : Sp12to4
    port map (
            O => \N__27982\,
            I => \N__27979\
        );

    \I__3902\ : Span12Mux_s9_h
    port map (
            O => \N__27979\,
            I => \N__27976\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__27976\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\
        );

    \I__3900\ : InMux
    port map (
            O => \N__27973\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__3899\ : InMux
    port map (
            O => \N__27970\,
            I => \N__27967\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__27967\,
            I => \N__27964\
        );

    \I__3897\ : Odrv12
    port map (
            O => \N__27964\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__3896\ : InMux
    port map (
            O => \N__27961\,
            I => \N__27958\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__27958\,
            I => \N__27955\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__27955\,
            I => \N__27952\
        );

    \I__3893\ : Sp12to4
    port map (
            O => \N__27952\,
            I => \N__27949\
        );

    \I__3892\ : Span12Mux_s9_h
    port map (
            O => \N__27949\,
            I => \N__27946\
        );

    \I__3891\ : Odrv12
    port map (
            O => \N__27946\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\
        );

    \I__3890\ : InMux
    port map (
            O => \N__27943\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__3889\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27934\
        );

    \I__3887\ : Sp12to4
    port map (
            O => \N__27934\,
            I => \N__27931\
        );

    \I__3886\ : Odrv12
    port map (
            O => \N__27931\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__3885\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27925\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__27925\,
            I => \N__27922\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__27922\,
            I => \N__27919\
        );

    \I__3882\ : Sp12to4
    port map (
            O => \N__27919\,
            I => \N__27916\
        );

    \I__3881\ : Span12Mux_s9_h
    port map (
            O => \N__27916\,
            I => \N__27913\
        );

    \I__3880\ : Odrv12
    port map (
            O => \N__27913\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\
        );

    \I__3879\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27906\
        );

    \I__3878\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27903\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__27906\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__27903\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\
        );

    \I__3875\ : InMux
    port map (
            O => \N__27898\,
            I => \bfn_9_14_0_\
        );

    \I__3874\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27892\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__27892\,
            I => \N__27889\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__27889\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\
        );

    \I__3871\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27882\
        );

    \I__3870\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27879\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__27882\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__27879\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\
        );

    \I__3867\ : InMux
    port map (
            O => \N__27874\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\
        );

    \I__3866\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27868\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__27862\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\
        );

    \I__3862\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27855\
        );

    \I__3861\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27852\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27847\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__27852\,
            I => \N__27847\
        );

    \I__3858\ : Span4Mux_v
    port map (
            O => \N__27847\,
            I => \N__27844\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__27844\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\
        );

    \I__3856\ : InMux
    port map (
            O => \N__27841\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\
        );

    \I__3855\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__27835\,
            I => \N__27831\
        );

    \I__3853\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27828\
        );

    \I__3852\ : Span4Mux_v
    port map (
            O => \N__27831\,
            I => \N__27825\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27822\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__27825\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__27822\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\
        );

    \I__3848\ : InMux
    port map (
            O => \N__27817\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\
        );

    \I__3847\ : InMux
    port map (
            O => \N__27814\,
            I => \N__27811\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__3845\ : Span4Mux_h
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__27805\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\
        );

    \I__3843\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27799\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27795\
        );

    \I__3841\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27792\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__27795\,
            I => \N__27789\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__27792\,
            I => \N__27786\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__27789\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__27786\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\
        );

    \I__3836\ : InMux
    port map (
            O => \N__27781\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\
        );

    \I__3835\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27774\
        );

    \I__3834\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27771\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__27774\,
            I => \N__27768\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__27771\,
            I => \N__27763\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__27768\,
            I => \N__27763\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__27763\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\
        );

    \I__3829\ : InMux
    port map (
            O => \N__27760\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\
        );

    \I__3828\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27754\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__27754\,
            I => \N__27751\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__27751\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\
        );

    \I__3825\ : InMux
    port map (
            O => \N__27748\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\
        );

    \I__3824\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27741\
        );

    \I__3823\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27738\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27735\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__27738\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__3820\ : Odrv12
    port map (
            O => \N__27735\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__3819\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27727\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__27727\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\
        );

    \I__3817\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27720\
        );

    \I__3816\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27717\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__27720\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__27717\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\
        );

    \I__3813\ : InMux
    port map (
            O => \N__27712\,
            I => \bfn_9_13_0_\
        );

    \I__3812\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27706\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__27706\,
            I => \N__27703\
        );

    \I__3810\ : Odrv12
    port map (
            O => \N__27703\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\
        );

    \I__3809\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27696\
        );

    \I__3808\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27693\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__27696\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__27693\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\
        );

    \I__3805\ : InMux
    port map (
            O => \N__27688\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\
        );

    \I__3804\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27682\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__27682\,
            I => \N__27679\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__27679\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\
        );

    \I__3801\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27672\
        );

    \I__3800\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27669\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__27672\,
            I => \N__27664\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__27669\,
            I => \N__27664\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__27664\,
            I => \N__27661\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__27661\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\
        );

    \I__3795\ : InMux
    port map (
            O => \N__27658\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\
        );

    \I__3794\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27648\
        );

    \I__3792\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27645\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__27648\,
            I => \N__27642\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27639\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__27642\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__27639\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\
        );

    \I__3787\ : InMux
    port map (
            O => \N__27634\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\
        );

    \I__3786\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27628\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__27628\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\
        );

    \I__3784\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27622\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27618\
        );

    \I__3782\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27615\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__27618\,
            I => \N__27612\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__27615\,
            I => \N__27609\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__27612\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__27609\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\
        );

    \I__3777\ : InMux
    port map (
            O => \N__27604\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\
        );

    \I__3776\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27597\
        );

    \I__3775\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27594\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__27597\,
            I => \N__27591\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27588\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__27591\,
            I => \N__27585\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__27588\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__27585\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\
        );

    \I__3769\ : InMux
    port map (
            O => \N__27580\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\
        );

    \I__3768\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27574\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27571\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__27571\,
            I => \N__27568\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__27568\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\
        );

    \I__3764\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27562\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__27562\,
            I => \N__27558\
        );

    \I__3762\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27555\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__27558\,
            I => \N__27550\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__27555\,
            I => \N__27550\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__27550\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\
        );

    \I__3758\ : InMux
    port map (
            O => \N__27547\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\
        );

    \I__3757\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27540\
        );

    \I__3756\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27537\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27534\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27529\
        );

    \I__3753\ : Span4Mux_h
    port map (
            O => \N__27534\,
            I => \N__27529\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__27529\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\
        );

    \I__3751\ : InMux
    port map (
            O => \N__27526\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\
        );

    \I__3750\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27520\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__27520\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\
        );

    \I__3748\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27514\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27510\
        );

    \I__3746\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27507\
        );

    \I__3745\ : Span4Mux_h
    port map (
            O => \N__27510\,
            I => \N__27504\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__27507\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__27504\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\
        );

    \I__3742\ : InMux
    port map (
            O => \N__27499\,
            I => \bfn_9_12_0_\
        );

    \I__3741\ : InMux
    port map (
            O => \N__27496\,
            I => \N__27493\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__27493\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\
        );

    \I__3739\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27486\
        );

    \I__3738\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27483\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__27486\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__27483\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\
        );

    \I__3735\ : InMux
    port map (
            O => \N__27478\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\
        );

    \I__3734\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27471\
        );

    \I__3733\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27468\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27463\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__27468\,
            I => \N__27463\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__27463\,
            I => \N__27460\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__27460\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\
        );

    \I__3728\ : InMux
    port map (
            O => \N__27457\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\
        );

    \I__3727\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27451\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__27451\,
            I => \N__27448\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__27448\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\
        );

    \I__3724\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27442\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27438\
        );

    \I__3722\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27435\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__27438\,
            I => \N__27432\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27429\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__27432\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__27429\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\
        );

    \I__3717\ : InMux
    port map (
            O => \N__27424\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\
        );

    \I__3716\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27414\
        );

    \I__3714\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27411\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__27414\,
            I => \N__27408\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27405\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__27408\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__27405\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\
        );

    \I__3709\ : InMux
    port map (
            O => \N__27400\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\
        );

    \I__3708\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27394\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__27394\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\
        );

    \I__3706\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27387\
        );

    \I__3705\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27384\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27381\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__27384\,
            I => \N__27376\
        );

    \I__3702\ : Span4Mux_h
    port map (
            O => \N__27381\,
            I => \N__27376\
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__27376\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\
        );

    \I__3700\ : InMux
    port map (
            O => \N__27373\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\
        );

    \I__3699\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__27367\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\
        );

    \I__3697\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__27361\,
            I => \N__27357\
        );

    \I__3695\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27354\
        );

    \I__3694\ : Span4Mux_h
    port map (
            O => \N__27357\,
            I => \N__27351\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__27354\,
            I => \N__27348\
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__27351\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__27348\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\
        );

    \I__3690\ : InMux
    port map (
            O => \N__27343\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\
        );

    \I__3689\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27337\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27334\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__27334\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\
        );

    \I__3686\ : InMux
    port map (
            O => \N__27331\,
            I => \N__27327\
        );

    \I__3685\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27324\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__27327\,
            I => \N__27321\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__27324\,
            I => \N__27316\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__27321\,
            I => \N__27316\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__27316\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\
        );

    \I__3680\ : InMux
    port map (
            O => \N__27313\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\
        );

    \I__3679\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27307\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__27307\,
            I => \N__27304\
        );

    \I__3677\ : Span4Mux_v
    port map (
            O => \N__27304\,
            I => \N__27300\
        );

    \I__3676\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27297\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__27300\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__27297\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__3673\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27289\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__27289\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__27286\,
            I => \N__27283\
        );

    \I__3670\ : InMux
    port map (
            O => \N__27283\,
            I => \N__27280\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__27280\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\
        );

    \I__3668\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27274\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__27274\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\
        );

    \I__3666\ : InMux
    port map (
            O => \N__27271\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\
        );

    \I__3665\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27265\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__27265\,
            I => \N__27261\
        );

    \I__3663\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27258\
        );

    \I__3662\ : Span4Mux_v
    port map (
            O => \N__27261\,
            I => \N__27255\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__27258\,
            I => \N__27252\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__27255\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__27252\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\
        );

    \I__3658\ : InMux
    port map (
            O => \N__27247\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\
        );

    \I__3657\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27241\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__27241\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\
        );

    \I__3655\ : InMux
    port map (
            O => \N__27238\,
            I => \N__27235\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__27235\,
            I => \N__27232\
        );

    \I__3653\ : Span4Mux_v
    port map (
            O => \N__27232\,
            I => \N__27228\
        );

    \I__3652\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27225\
        );

    \I__3651\ : Span4Mux_v
    port map (
            O => \N__27228\,
            I => \N__27220\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__27225\,
            I => \N__27220\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__27220\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\
        );

    \I__3648\ : InMux
    port map (
            O => \N__27217\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\
        );

    \I__3647\ : InMux
    port map (
            O => \N__27214\,
            I => \N__27210\
        );

    \I__3646\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27207\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__27210\,
            I => \N__27204\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27201\
        );

    \I__3643\ : Span4Mux_h
    port map (
            O => \N__27204\,
            I => \N__27198\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__27201\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__27198\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\
        );

    \I__3640\ : InMux
    port map (
            O => \N__27193\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\
        );

    \I__3639\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__27184\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\
        );

    \I__3636\ : InMux
    port map (
            O => \N__27181\,
            I => \N__27178\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__27178\,
            I => \N__27174\
        );

    \I__3634\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27171\
        );

    \I__3633\ : Span4Mux_h
    port map (
            O => \N__27174\,
            I => \N__27168\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27165\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__27168\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__27165\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\
        );

    \I__3629\ : InMux
    port map (
            O => \N__27160\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\
        );

    \I__3628\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27153\
        );

    \I__3627\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27150\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__27153\,
            I => \N__27145\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27145\
        );

    \I__3624\ : Span4Mux_h
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__27142\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\
        );

    \I__3622\ : InMux
    port map (
            O => \N__27139\,
            I => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\
        );

    \I__3621\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27130\
        );

    \I__3620\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27130\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__27130\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__3618\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27123\
        );

    \I__3617\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27120\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__27123\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__27120\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__3614\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27112\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__27112\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__27109\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\
        );

    \I__3611\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27102\
        );

    \I__3610\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27099\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__27102\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__27099\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__3607\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27091\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27087\
        );

    \I__3605\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27084\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__27087\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__27084\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__3602\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27076\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__27076\,
            I => \N__27072\
        );

    \I__3600\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27069\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__27072\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__27069\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__3597\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__27061\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__3595\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27055\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__27055\,
            I => \N__27051\
        );

    \I__3593\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27048\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__27051\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__27048\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__3590\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27040\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__27040\,
            I => \N__27037\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__27037\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__27034\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5_cascade_\
        );

    \I__3586\ : InMux
    port map (
            O => \N__27031\,
            I => \N__27027\
        );

    \I__3585\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27024\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__27027\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__27024\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__27019\,
            I => \N__27015\
        );

    \I__3581\ : InMux
    port map (
            O => \N__27018\,
            I => \N__27012\
        );

    \I__3580\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27009\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__27012\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__27009\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__3577\ : InMux
    port map (
            O => \N__27004\,
            I => \N__27001\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__27001\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__3575\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26994\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__26997\,
            I => \N__26991\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__26994\,
            I => \N__26988\
        );

    \I__3572\ : InMux
    port map (
            O => \N__26991\,
            I => \N__26985\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__26988\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__26985\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__26980\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\
        );

    \I__3568\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26971\
        );

    \I__3567\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26971\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__26971\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__3565\ : InMux
    port map (
            O => \N__26968\,
            I => \N__26964\
        );

    \I__3564\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26961\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__26964\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__26961\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__3561\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26949\
        );

    \I__3559\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26946\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__26949\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__26946\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__3556\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26937\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__26940\,
            I => \N__26934\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26931\
        );

    \I__3553\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26928\
        );

    \I__3552\ : Odrv12
    port map (
            O => \N__26931\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__26928\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__3550\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26917\
        );

    \I__3549\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26917\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__26917\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__3547\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26907\
        );

    \I__3545\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26904\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__26907\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__26904\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__26899\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\
        );

    \I__3541\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26886\
        );

    \I__3540\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26886\
        );

    \I__3539\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26886\
        );

    \I__3538\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26883\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__26886\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__26883\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__26878\,
            I => \N__26874\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__26877\,
            I => \N__26871\
        );

    \I__3533\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26862\
        );

    \I__3532\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26862\
        );

    \I__3531\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26862\
        );

    \I__3530\ : InMux
    port map (
            O => \N__26869\,
            I => \N__26859\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__26862\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__26859\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__3527\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26851\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__26851\,
            I => \phase_controller_inst2.start_timer_tr_0_sqmuxa\
        );

    \I__3525\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26845\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__26845\,
            I => \N__26842\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__26842\,
            I => \N__26839\
        );

    \I__3522\ : Sp12to4
    port map (
            O => \N__26839\,
            I => \N__26836\
        );

    \I__3521\ : Span12Mux_h
    port map (
            O => \N__26836\,
            I => \N__26833\
        );

    \I__3520\ : Odrv12
    port map (
            O => \N__26833\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__3519\ : InMux
    port map (
            O => \N__26830\,
            I => \bfn_8_22_0_\
        );

    \I__3518\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26824\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__26824\,
            I => \N__26821\
        );

    \I__3516\ : Span12Mux_v
    port map (
            O => \N__26821\,
            I => \N__26818\
        );

    \I__3515\ : Span12Mux_h
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__3514\ : Odrv12
    port map (
            O => \N__26815\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__3513\ : InMux
    port map (
            O => \N__26812\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__3512\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26806\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__26806\,
            I => \N__26803\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__26803\,
            I => \N__26800\
        );

    \I__3509\ : Sp12to4
    port map (
            O => \N__26800\,
            I => \N__26797\
        );

    \I__3508\ : Span12Mux_h
    port map (
            O => \N__26797\,
            I => \N__26794\
        );

    \I__3507\ : Odrv12
    port map (
            O => \N__26794\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__3506\ : InMux
    port map (
            O => \N__26791\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__3505\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26785\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__26785\,
            I => \N__26782\
        );

    \I__3503\ : Span4Mux_v
    port map (
            O => \N__26782\,
            I => \N__26779\
        );

    \I__3502\ : Sp12to4
    port map (
            O => \N__26779\,
            I => \N__26776\
        );

    \I__3501\ : Span12Mux_h
    port map (
            O => \N__26776\,
            I => \N__26773\
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__26773\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__3499\ : InMux
    port map (
            O => \N__26770\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__3498\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26764\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__26764\,
            I => \N__26761\
        );

    \I__3496\ : Span4Mux_v
    port map (
            O => \N__26761\,
            I => \N__26758\
        );

    \I__3495\ : Sp12to4
    port map (
            O => \N__26758\,
            I => \N__26755\
        );

    \I__3494\ : Span12Mux_h
    port map (
            O => \N__26755\,
            I => \N__26752\
        );

    \I__3493\ : Odrv12
    port map (
            O => \N__26752\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__3492\ : InMux
    port map (
            O => \N__26749\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__3491\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26743\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__26743\,
            I => \N__26740\
        );

    \I__3489\ : Span4Mux_v
    port map (
            O => \N__26740\,
            I => \N__26737\
        );

    \I__3488\ : Sp12to4
    port map (
            O => \N__26737\,
            I => \N__26734\
        );

    \I__3487\ : Span12Mux_h
    port map (
            O => \N__26734\,
            I => \N__26731\
        );

    \I__3486\ : Odrv12
    port map (
            O => \N__26731\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26728\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__3484\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26722\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__26722\,
            I => \N__26719\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__26719\,
            I => \N__26716\
        );

    \I__3481\ : Sp12to4
    port map (
            O => \N__26716\,
            I => \N__26713\
        );

    \I__3480\ : Span12Mux_h
    port map (
            O => \N__26713\,
            I => \N__26710\
        );

    \I__3479\ : Odrv12
    port map (
            O => \N__26710\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__3478\ : InMux
    port map (
            O => \N__26707\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__3477\ : InMux
    port map (
            O => \N__26704\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__3476\ : InMux
    port map (
            O => \N__26701\,
            I => \N__26698\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__26698\,
            I => \N__26695\
        );

    \I__3474\ : Span4Mux_v
    port map (
            O => \N__26695\,
            I => \N__26692\
        );

    \I__3473\ : Sp12to4
    port map (
            O => \N__26692\,
            I => \N__26689\
        );

    \I__3472\ : Span12Mux_h
    port map (
            O => \N__26689\,
            I => \N__26686\
        );

    \I__3471\ : Odrv12
    port map (
            O => \N__26686\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__26683\,
            I => \N__26680\
        );

    \I__3469\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26674\
        );

    \I__3467\ : Span4Mux_v
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__3466\ : Sp12to4
    port map (
            O => \N__26671\,
            I => \N__26668\
        );

    \I__3465\ : Span12Mux_v
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__3464\ : Odrv12
    port map (
            O => \N__26665\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__3463\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26659\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26656\
        );

    \I__3461\ : Span12Mux_v
    port map (
            O => \N__26656\,
            I => \N__26653\
        );

    \I__3460\ : Span12Mux_h
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__3459\ : Odrv12
    port map (
            O => \N__26650\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__26647\,
            I => \N__26644\
        );

    \I__3457\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26641\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__26641\,
            I => \N__26638\
        );

    \I__3455\ : Span12Mux_s11_v
    port map (
            O => \N__26638\,
            I => \N__26635\
        );

    \I__3454\ : Span12Mux_v
    port map (
            O => \N__26635\,
            I => \N__26632\
        );

    \I__3453\ : Odrv12
    port map (
            O => \N__26632\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__3452\ : InMux
    port map (
            O => \N__26629\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__3451\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26620\
        );

    \I__3449\ : Span12Mux_h
    port map (
            O => \N__26620\,
            I => \N__26617\
        );

    \I__3448\ : Span12Mux_h
    port map (
            O => \N__26617\,
            I => \N__26614\
        );

    \I__3447\ : Odrv12
    port map (
            O => \N__26614\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__3445\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26605\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__26605\,
            I => \N__26602\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__26602\,
            I => \N__26599\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__26599\,
            I => \N__26596\
        );

    \I__3441\ : Span4Mux_h
    port map (
            O => \N__26596\,
            I => \N__26593\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__26593\,
            I => \N__26590\
        );

    \I__3439\ : Span4Mux_v
    port map (
            O => \N__26590\,
            I => \N__26587\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__26587\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__3437\ : InMux
    port map (
            O => \N__26584\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__3436\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26575\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__26575\,
            I => \N__26572\
        );

    \I__3433\ : Sp12to4
    port map (
            O => \N__26572\,
            I => \N__26569\
        );

    \I__3432\ : Span12Mux_h
    port map (
            O => \N__26569\,
            I => \N__26566\
        );

    \I__3431\ : Odrv12
    port map (
            O => \N__26566\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__26563\,
            I => \N__26560\
        );

    \I__3429\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26557\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__26557\,
            I => \N__26554\
        );

    \I__3427\ : Span12Mux_h
    port map (
            O => \N__26554\,
            I => \N__26551\
        );

    \I__3426\ : Span12Mux_v
    port map (
            O => \N__26551\,
            I => \N__26548\
        );

    \I__3425\ : Odrv12
    port map (
            O => \N__26548\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__3424\ : InMux
    port map (
            O => \N__26545\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__3423\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__26539\,
            I => \N__26536\
        );

    \I__3421\ : Span4Mux_v
    port map (
            O => \N__26536\,
            I => \N__26533\
        );

    \I__3420\ : Sp12to4
    port map (
            O => \N__26533\,
            I => \N__26530\
        );

    \I__3419\ : Span12Mux_h
    port map (
            O => \N__26530\,
            I => \N__26527\
        );

    \I__3418\ : Odrv12
    port map (
            O => \N__26527\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__3417\ : InMux
    port map (
            O => \N__26524\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26518\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__26518\,
            I => \N__26515\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__26515\,
            I => \N__26512\
        );

    \I__3413\ : Sp12to4
    port map (
            O => \N__26512\,
            I => \N__26509\
        );

    \I__3412\ : Span12Mux_h
    port map (
            O => \N__26509\,
            I => \N__26506\
        );

    \I__3411\ : Odrv12
    port map (
            O => \N__26506\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__3410\ : InMux
    port map (
            O => \N__26503\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__3409\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26497\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__26497\,
            I => \N__26494\
        );

    \I__3407\ : Span4Mux_v
    port map (
            O => \N__26494\,
            I => \N__26491\
        );

    \I__3406\ : Sp12to4
    port map (
            O => \N__26491\,
            I => \N__26488\
        );

    \I__3405\ : Span12Mux_h
    port map (
            O => \N__26488\,
            I => \N__26485\
        );

    \I__3404\ : Odrv12
    port map (
            O => \N__26485\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__3403\ : InMux
    port map (
            O => \N__26482\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__3402\ : InMux
    port map (
            O => \N__26479\,
            I => \N__26476\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__26476\,
            I => \N__26473\
        );

    \I__3400\ : Span4Mux_v
    port map (
            O => \N__26473\,
            I => \N__26470\
        );

    \I__3399\ : Sp12to4
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__3398\ : Span12Mux_h
    port map (
            O => \N__26467\,
            I => \N__26464\
        );

    \I__3397\ : Odrv12
    port map (
            O => \N__26464\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__3396\ : InMux
    port map (
            O => \N__26461\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__3395\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26452\
        );

    \I__3394\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26452\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26448\
        );

    \I__3392\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26445\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__26448\,
            I => \N__26442\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__26445\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_24\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__26442\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_24\
        );

    \I__3388\ : InMux
    port map (
            O => \N__26437\,
            I => \bfn_8_20_0_\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__26434\,
            I => \N__26430\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__26433\,
            I => \N__26427\
        );

    \I__3385\ : InMux
    port map (
            O => \N__26430\,
            I => \N__26422\
        );

    \I__3384\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26422\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__26422\,
            I => \N__26418\
        );

    \I__3382\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26415\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__26418\,
            I => \N__26412\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__26415\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_25\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__26412\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_25\
        );

    \I__3378\ : InMux
    port map (
            O => \N__26407\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_24\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__26404\,
            I => \N__26400\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__26403\,
            I => \N__26397\
        );

    \I__3375\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26392\
        );

    \I__3374\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26392\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__26392\,
            I => \N__26388\
        );

    \I__3372\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26385\
        );

    \I__3371\ : Span4Mux_h
    port map (
            O => \N__26388\,
            I => \N__26382\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__26385\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_26\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__26382\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_26\
        );

    \I__3368\ : InMux
    port map (
            O => \N__26377\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_25\
        );

    \I__3367\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26368\
        );

    \I__3366\ : InMux
    port map (
            O => \N__26373\,
            I => \N__26368\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__26368\,
            I => \N__26364\
        );

    \I__3364\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26361\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__26364\,
            I => \N__26358\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__26361\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__26358\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_27\
        );

    \I__3360\ : InMux
    port map (
            O => \N__26353\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_26\
        );

    \I__3359\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26345\
        );

    \I__3358\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26342\
        );

    \I__3357\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26339\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__26345\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__26342\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__26339\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_28\
        );

    \I__3353\ : InMux
    port map (
            O => \N__26332\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_27\
        );

    \I__3352\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26324\
        );

    \I__3351\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26319\
        );

    \I__3350\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26319\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__26324\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__26319\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_29\
        );

    \I__3347\ : InMux
    port map (
            O => \N__26314\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_28\
        );

    \I__3346\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26306\
        );

    \I__3345\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26301\
        );

    \I__3344\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26301\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__26306\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__26301\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_30\
        );

    \I__3341\ : InMux
    port map (
            O => \N__26296\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_29\
        );

    \I__3340\ : InMux
    port map (
            O => \N__26293\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_30\
        );

    \I__3339\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26285\
        );

    \I__3338\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26282\
        );

    \I__3337\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26279\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__26285\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__26282\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__26279\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_31\
        );

    \I__3333\ : CEMux
    port map (
            O => \N__26272\,
            I => \N__26260\
        );

    \I__3332\ : CEMux
    port map (
            O => \N__26271\,
            I => \N__26260\
        );

    \I__3331\ : CEMux
    port map (
            O => \N__26270\,
            I => \N__26260\
        );

    \I__3330\ : CEMux
    port map (
            O => \N__26269\,
            I => \N__26260\
        );

    \I__3329\ : GlobalMux
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__3328\ : gio2CtrlBuf
    port map (
            O => \N__26257\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0_g\
        );

    \I__3327\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26250\
        );

    \I__3326\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26247\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__26250\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_15\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__26247\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_15\
        );

    \I__3323\ : InMux
    port map (
            O => \N__26242\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_14\
        );

    \I__3322\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26233\
        );

    \I__3321\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26233\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__26233\,
            I => \N__26229\
        );

    \I__3319\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26226\
        );

    \I__3318\ : Span4Mux_v
    port map (
            O => \N__26229\,
            I => \N__26223\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__26226\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_16\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__26223\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_16\
        );

    \I__3315\ : InMux
    port map (
            O => \N__26218\,
            I => \bfn_8_19_0_\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \N__26211\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__26214\,
            I => \N__26208\
        );

    \I__3312\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26203\
        );

    \I__3311\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26203\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26199\
        );

    \I__3309\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26196\
        );

    \I__3308\ : Span4Mux_v
    port map (
            O => \N__26199\,
            I => \N__26193\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__26196\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_17\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__26193\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_17\
        );

    \I__3305\ : InMux
    port map (
            O => \N__26188\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_16\
        );

    \I__3304\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26179\
        );

    \I__3303\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26179\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__26179\,
            I => \N__26175\
        );

    \I__3301\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26172\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__26175\,
            I => \N__26169\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__26172\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_18\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__26169\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_18\
        );

    \I__3297\ : InMux
    port map (
            O => \N__26164\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_17\
        );

    \I__3296\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26155\
        );

    \I__3295\ : InMux
    port map (
            O => \N__26160\,
            I => \N__26155\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__26155\,
            I => \N__26151\
        );

    \I__3293\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26148\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__26151\,
            I => \N__26145\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__26148\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_19\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__26145\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_19\
        );

    \I__3289\ : InMux
    port map (
            O => \N__26140\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_18\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__26137\,
            I => \N__26133\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__26136\,
            I => \N__26130\
        );

    \I__3286\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26124\
        );

    \I__3285\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26124\
        );

    \I__3284\ : InMux
    port map (
            O => \N__26129\,
            I => \N__26121\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__26124\,
            I => \N__26118\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__26121\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_20\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__26118\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_20\
        );

    \I__3280\ : InMux
    port map (
            O => \N__26113\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_19\
        );

    \I__3279\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26103\
        );

    \I__3278\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26103\
        );

    \I__3277\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26100\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__26103\,
            I => \N__26097\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__26100\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_21\
        );

    \I__3274\ : Odrv4
    port map (
            O => \N__26097\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_21\
        );

    \I__3273\ : InMux
    port map (
            O => \N__26092\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_20\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__26089\,
            I => \N__26085\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__26088\,
            I => \N__26082\
        );

    \I__3270\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26077\
        );

    \I__3269\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26077\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__26077\,
            I => \N__26073\
        );

    \I__3267\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26070\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__26073\,
            I => \N__26067\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__26070\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_22\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__26067\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_22\
        );

    \I__3263\ : InMux
    port map (
            O => \N__26062\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_21\
        );

    \I__3262\ : InMux
    port map (
            O => \N__26059\,
            I => \N__26053\
        );

    \I__3261\ : InMux
    port map (
            O => \N__26058\,
            I => \N__26053\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__26053\,
            I => \N__26049\
        );

    \I__3259\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26046\
        );

    \I__3258\ : Span4Mux_h
    port map (
            O => \N__26049\,
            I => \N__26043\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__26046\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_23\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__26043\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_23\
        );

    \I__3255\ : InMux
    port map (
            O => \N__26038\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_22\
        );

    \I__3254\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26031\
        );

    \I__3253\ : InMux
    port map (
            O => \N__26034\,
            I => \N__26028\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__26031\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_7\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__26028\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_7\
        );

    \I__3250\ : InMux
    port map (
            O => \N__26023\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_6\
        );

    \I__3249\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26016\
        );

    \I__3248\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26013\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__26016\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_8\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__26013\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_8\
        );

    \I__3245\ : InMux
    port map (
            O => \N__26008\,
            I => \bfn_8_18_0_\
        );

    \I__3244\ : InMux
    port map (
            O => \N__26005\,
            I => \N__26001\
        );

    \I__3243\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25998\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__26001\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_9\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__25998\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_9\
        );

    \I__3240\ : InMux
    port map (
            O => \N__25993\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_8\
        );

    \I__3239\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25986\
        );

    \I__3238\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25983\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__25986\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_10\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__25983\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_10\
        );

    \I__3235\ : InMux
    port map (
            O => \N__25978\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_9\
        );

    \I__3234\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25971\
        );

    \I__3233\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25968\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__25971\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_11\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__25968\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_11\
        );

    \I__3230\ : InMux
    port map (
            O => \N__25963\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_10\
        );

    \I__3229\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25956\
        );

    \I__3228\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25953\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__25956\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_12\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__25953\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_12\
        );

    \I__3225\ : InMux
    port map (
            O => \N__25948\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_11\
        );

    \I__3224\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25941\
        );

    \I__3223\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25938\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__25941\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_13\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__25938\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_13\
        );

    \I__3220\ : InMux
    port map (
            O => \N__25933\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_12\
        );

    \I__3219\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25926\
        );

    \I__3218\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25923\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__25926\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_14\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__25923\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_14\
        );

    \I__3215\ : InMux
    port map (
            O => \N__25918\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_13\
        );

    \I__3214\ : InMux
    port map (
            O => \N__25915\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__25912\,
            I => \N__25908\
        );

    \I__3212\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25905\
        );

    \I__3211\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25902\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25897\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25897\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__25897\,
            I => \phase_controller_inst2.stoper_tr.counter\
        );

    \I__3207\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25890\
        );

    \I__3206\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25887\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__25890\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_0\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__25887\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_0\
        );

    \I__3203\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25878\
        );

    \I__3202\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25875\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__25878\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_1\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25875\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_1\
        );

    \I__3199\ : InMux
    port map (
            O => \N__25870\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_0\
        );

    \I__3198\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25863\
        );

    \I__3197\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25860\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__25863\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_2\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__25860\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_2\
        );

    \I__3194\ : InMux
    port map (
            O => \N__25855\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_1\
        );

    \I__3193\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25848\
        );

    \I__3192\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25845\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__25848\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_3\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__25845\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_3\
        );

    \I__3189\ : InMux
    port map (
            O => \N__25840\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_2\
        );

    \I__3188\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25833\
        );

    \I__3187\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25830\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__25833\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_4\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__25830\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_4\
        );

    \I__3184\ : InMux
    port map (
            O => \N__25825\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_3\
        );

    \I__3183\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25818\
        );

    \I__3182\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25815\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__25818\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_5\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__25815\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_5\
        );

    \I__3179\ : InMux
    port map (
            O => \N__25810\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_4\
        );

    \I__3178\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25803\
        );

    \I__3177\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25800\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__25803\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_6\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__25800\,
            I => \phase_controller_inst2.stoper_tr.counterZ0Z_6\
        );

    \I__3174\ : InMux
    port map (
            O => \N__25795\,
            I => \phase_controller_inst2.stoper_tr.counter_cry_5\
        );

    \I__3173\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25789\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25785\
        );

    \I__3171\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25782\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__25785\,
            I => \N__25777\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__25782\,
            I => \N__25777\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__25777\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_19
        );

    \I__3167\ : InMux
    port map (
            O => \N__25774\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\
        );

    \I__3166\ : InMux
    port map (
            O => \N__25771\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\
        );

    \I__3165\ : InMux
    port map (
            O => \N__25768\,
            I => \N__25765\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__25762\,
            I => \N__25758\
        );

    \I__3162\ : InMux
    port map (
            O => \N__25761\,
            I => \N__25755\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__25758\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_21
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__25755\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_21
        );

    \I__3159\ : InMux
    port map (
            O => \N__25750\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\
        );

    \I__3158\ : InMux
    port map (
            O => \N__25747\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\
        );

    \I__3157\ : InMux
    port map (
            O => \N__25744\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\
        );

    \I__3156\ : InMux
    port map (
            O => \N__25741\,
            I => \bfn_8_16_0_\
        );

    \I__3155\ : InMux
    port map (
            O => \N__25738\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\
        );

    \I__3154\ : InMux
    port map (
            O => \N__25735\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\
        );

    \I__3153\ : InMux
    port map (
            O => \N__25732\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\
        );

    \I__3152\ : InMux
    port map (
            O => \N__25729\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\
        );

    \I__3151\ : InMux
    port map (
            O => \N__25726\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\
        );

    \I__3150\ : InMux
    port map (
            O => \N__25723\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\
        );

    \I__3149\ : InMux
    port map (
            O => \N__25720\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\
        );

    \I__3148\ : InMux
    port map (
            O => \N__25717\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\
        );

    \I__3147\ : InMux
    port map (
            O => \N__25714\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\
        );

    \I__3146\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25708\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__25705\,
            I => \N__25701\
        );

    \I__3143\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25698\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__25701\,
            I => \N__25695\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__25698\,
            I => \N__25692\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__25695\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_16
        );

    \I__3139\ : Odrv12
    port map (
            O => \N__25692\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_16
        );

    \I__3138\ : InMux
    port map (
            O => \N__25687\,
            I => \bfn_8_15_0_\
        );

    \I__3137\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25681\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__25681\,
            I => \N__25677\
        );

    \I__3135\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25674\
        );

    \I__3134\ : Span4Mux_v
    port map (
            O => \N__25677\,
            I => \N__25671\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__25674\,
            I => \N__25668\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__25671\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_17
        );

    \I__3131\ : Odrv12
    port map (
            O => \N__25668\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_17
        );

    \I__3130\ : InMux
    port map (
            O => \N__25663\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\
        );

    \I__3129\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25653\
        );

    \I__3127\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25650\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__25653\,
            I => \N__25645\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__25650\,
            I => \N__25645\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__25645\,
            I => phase_controller_inst1_stoper_tr_target_ticks_1_i_18
        );

    \I__3123\ : InMux
    port map (
            O => \N__25642\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\
        );

    \I__3122\ : InMux
    port map (
            O => \N__25639\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\
        );

    \I__3121\ : InMux
    port map (
            O => \N__25636\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\
        );

    \I__3120\ : InMux
    port map (
            O => \N__25633\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\
        );

    \I__3119\ : InMux
    port map (
            O => \N__25630\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\
        );

    \I__3118\ : InMux
    port map (
            O => \N__25627\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\
        );

    \I__3117\ : InMux
    port map (
            O => \N__25624\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\
        );

    \I__3116\ : InMux
    port map (
            O => \N__25621\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\
        );

    \I__3115\ : InMux
    port map (
            O => \N__25618\,
            I => \bfn_8_14_0_\
        );

    \I__3114\ : InMux
    port map (
            O => \N__25615\,
            I => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\
        );

    \I__3113\ : InMux
    port map (
            O => \N__25612\,
            I => \N__25608\
        );

    \I__3112\ : InMux
    port map (
            O => \N__25611\,
            I => \N__25605\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__25608\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__25605\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__3109\ : InMux
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__25597\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__25594\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\
        );

    \I__3106\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25587\
        );

    \I__3105\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25584\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__25587\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__25584\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3102\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25576\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__25576\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__25573\,
            I => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\
        );

    \I__3099\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25566\
        );

    \I__3098\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25563\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__25566\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__25563\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__3095\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25555\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__25555\,
            I => \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__25552\,
            I => \N__25549\
        );

    \I__3092\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25544\
        );

    \I__3091\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25541\
        );

    \I__3090\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25538\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__25544\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__25541\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__25538\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__3086\ : InMux
    port map (
            O => \N__25531\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__3084\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25520\
        );

    \I__3083\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25517\
        );

    \I__3082\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25514\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__25520\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__25517\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__25514\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__3078\ : InMux
    port map (
            O => \N__25507\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__25504\,
            I => \N__25501\
        );

    \I__3076\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25496\
        );

    \I__3075\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25493\
        );

    \I__3074\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25490\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__25496\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__25493\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__25490\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__3070\ : InMux
    port map (
            O => \N__25483\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__25480\,
            I => \N__25477\
        );

    \I__3068\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25472\
        );

    \I__3067\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25469\
        );

    \I__3066\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25466\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__25472\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__25469\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__25466\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__3062\ : InMux
    port map (
            O => \N__25459\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__25456\,
            I => \N__25453\
        );

    \I__3060\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25448\
        );

    \I__3059\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25445\
        );

    \I__3058\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25442\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__25448\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__25445\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__25442\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__3054\ : InMux
    port map (
            O => \N__25435\,
            I => \bfn_8_11_0_\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__25432\,
            I => \N__25429\
        );

    \I__3052\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25424\
        );

    \I__3051\ : InMux
    port map (
            O => \N__25428\,
            I => \N__25421\
        );

    \I__3050\ : InMux
    port map (
            O => \N__25427\,
            I => \N__25418\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__25424\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__25421\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__25418\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__3046\ : InMux
    port map (
            O => \N__25411\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__3045\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25404\
        );

    \I__3044\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25401\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__25404\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__25401\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__3040\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25388\
        );

    \I__3039\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25385\
        );

    \I__3038\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25382\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__25388\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__25385\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__25382\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__3034\ : InMux
    port map (
            O => \N__25375\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__3033\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25368\
        );

    \I__3032\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25365\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__25368\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__25365\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__25360\,
            I => \N__25357\
        );

    \I__3028\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25352\
        );

    \I__3027\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25349\
        );

    \I__3026\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25346\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__25352\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__25349\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__25346\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__3022\ : InMux
    port map (
            O => \N__25339\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__3021\ : InMux
    port map (
            O => \N__25336\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__25333\,
            I => \N__25330\
        );

    \I__3019\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25325\
        );

    \I__3018\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25322\
        );

    \I__3017\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25319\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__25325\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__25322\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__25319\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__3013\ : InMux
    port map (
            O => \N__25312\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__25309\,
            I => \N__25306\
        );

    \I__3011\ : InMux
    port map (
            O => \N__25306\,
            I => \N__25301\
        );

    \I__3010\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25298\
        );

    \I__3009\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25295\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__25301\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__25298\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__25295\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__3005\ : InMux
    port map (
            O => \N__25288\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__25285\,
            I => \N__25282\
        );

    \I__3003\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25277\
        );

    \I__3002\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25274\
        );

    \I__3001\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25271\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__25277\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__25274\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__25271\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__2997\ : InMux
    port map (
            O => \N__25264\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__25261\,
            I => \N__25258\
        );

    \I__2995\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25253\
        );

    \I__2994\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25250\
        );

    \I__2993\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25247\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__25253\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__25250\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__25247\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__2989\ : InMux
    port map (
            O => \N__25240\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__25237\,
            I => \N__25234\
        );

    \I__2987\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25229\
        );

    \I__2986\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25226\
        );

    \I__2985\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25223\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__25229\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__25226\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__25223\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__2981\ : InMux
    port map (
            O => \N__25216\,
            I => \bfn_8_10_0_\
        );

    \I__2980\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25208\
        );

    \I__2979\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25205\
        );

    \I__2978\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25202\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__25208\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__25205\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__25202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__2974\ : InMux
    port map (
            O => \N__25195\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__25192\,
            I => \N__25189\
        );

    \I__2972\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25184\
        );

    \I__2971\ : InMux
    port map (
            O => \N__25188\,
            I => \N__25181\
        );

    \I__2970\ : InMux
    port map (
            O => \N__25187\,
            I => \N__25178\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__25184\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__25181\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__25178\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__2966\ : InMux
    port map (
            O => \N__25171\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__25168\,
            I => \N__25163\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__25167\,
            I => \N__25160\
        );

    \I__2963\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25157\
        );

    \I__2962\ : InMux
    port map (
            O => \N__25163\,
            I => \N__25152\
        );

    \I__2961\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25152\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__25157\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__25152\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__2958\ : InMux
    port map (
            O => \N__25147\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__2957\ : InMux
    port map (
            O => \N__25144\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__25141\,
            I => \N__25136\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__25140\,
            I => \N__25133\
        );

    \I__2954\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25130\
        );

    \I__2953\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25125\
        );

    \I__2952\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25125\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__25130\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__25125\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__2949\ : InMux
    port map (
            O => \N__25120\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__25117\,
            I => \N__25114\
        );

    \I__2947\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25109\
        );

    \I__2946\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25106\
        );

    \I__2945\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25103\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__25109\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__25106\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__25103\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__2941\ : InMux
    port map (
            O => \N__25096\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__25093\,
            I => \N__25090\
        );

    \I__2939\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25085\
        );

    \I__2938\ : InMux
    port map (
            O => \N__25089\,
            I => \N__25082\
        );

    \I__2937\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25079\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__25085\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__25082\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__25079\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__2933\ : InMux
    port map (
            O => \N__25072\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__25069\,
            I => \N__25066\
        );

    \I__2931\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25061\
        );

    \I__2930\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25058\
        );

    \I__2929\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25055\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__25061\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__25058\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__25055\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__2925\ : InMux
    port map (
            O => \N__25048\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__25045\,
            I => \N__25042\
        );

    \I__2923\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25037\
        );

    \I__2922\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25034\
        );

    \I__2921\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25031\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__25037\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__25034\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__25031\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__2917\ : InMux
    port map (
            O => \N__25024\,
            I => \bfn_8_9_0_\
        );

    \I__2916\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25016\
        );

    \I__2915\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25013\
        );

    \I__2914\ : InMux
    port map (
            O => \N__25019\,
            I => \N__25010\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__25016\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__25013\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__25010\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__2910\ : InMux
    port map (
            O => \N__25003\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__2908\ : InMux
    port map (
            O => \N__24997\,
            I => \N__24992\
        );

    \I__2907\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24989\
        );

    \I__2906\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24986\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__24992\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__24989\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__24986\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__2902\ : InMux
    port map (
            O => \N__24979\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__24976\,
            I => \N__24971\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__24975\,
            I => \N__24968\
        );

    \I__2899\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24965\
        );

    \I__2898\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24960\
        );

    \I__2897\ : InMux
    port map (
            O => \N__24968\,
            I => \N__24960\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__24965\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__24960\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__2894\ : InMux
    port map (
            O => \N__24955\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__2893\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24949\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__24949\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt30\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__2890\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__24940\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\
        );

    \I__2888\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__24934\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt28\
        );

    \I__2886\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24928\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24925\
        );

    \I__2884\ : Glb2LocalMux
    port map (
            O => \N__24925\,
            I => \N__24922\
        );

    \I__2883\ : GlobalMux
    port map (
            O => \N__24922\,
            I => clk_12mhz
        );

    \I__2882\ : IoInMux
    port map (
            O => \N__24919\,
            I => \N__24916\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__24916\,
            I => \N__24913\
        );

    \I__2880\ : Span4Mux_s0_v
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__2879\ : Odrv4
    port map (
            O => \N__24910\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2878\ : InMux
    port map (
            O => \N__24907\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__2877\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24899\
        );

    \I__2876\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24894\
        );

    \I__2875\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24894\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__24899\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__24894\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__2872\ : InMux
    port map (
            O => \N__24889\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__2870\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24878\
        );

    \I__2869\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24875\
        );

    \I__2868\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24872\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__24878\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__24875\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__24872\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__2864\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24862\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__24862\,
            I => \N__24859\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__24859\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__24856\,
            I => \N__24853\
        );

    \I__2860\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24850\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24847\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__24847\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt20\
        );

    \I__2857\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24841\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__24841\,
            I => \N__24838\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__24835\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__24832\,
            I => \N__24829\
        );

    \I__2852\ : InMux
    port map (
            O => \N__24829\,
            I => \N__24826\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24823\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__24823\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt22\
        );

    \I__2849\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24817\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__24817\,
            I => \N__24814\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__24814\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__24811\,
            I => \N__24808\
        );

    \I__2845\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24805\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__24805\,
            I => \N__24802\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__24802\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt24\
        );

    \I__2842\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24796\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__24796\,
            I => \N__24793\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__24793\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__2838\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24784\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__24784\,
            I => \N__24781\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__24781\,
            I => \N__24778\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__24778\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt26\
        );

    \I__2834\ : InMux
    port map (
            O => \N__24775\,
            I => \bfn_7_20_0_\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \N__24769\
        );

    \I__2832\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__24766\,
            I => \N__24763\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__24763\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\
        );

    \I__2829\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24757\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24754\
        );

    \I__2827\ : Odrv12
    port map (
            O => \N__24754\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__24751\,
            I => \N__24748\
        );

    \I__2825\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24745\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__24745\,
            I => \phase_controller_inst2.stoper_tr.counter_i_10\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__2822\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24736\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24733\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__24733\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\
        );

    \I__2819\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24727\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__24727\,
            I => \phase_controller_inst2.stoper_tr.counter_i_11\
        );

    \I__2817\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24721\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__24721\,
            I => \N__24718\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__24718\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__24715\,
            I => \N__24712\
        );

    \I__2813\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24709\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__24709\,
            I => \phase_controller_inst2.stoper_tr.counter_i_12\
        );

    \I__2811\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24703\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__24703\,
            I => \N__24700\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__24700\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__24697\,
            I => \N__24694\
        );

    \I__2807\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__24691\,
            I => \N__24688\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__24688\,
            I => \phase_controller_inst2.stoper_tr.counter_i_13\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__24685\,
            I => \N__24682\
        );

    \I__2803\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24679\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__24679\,
            I => \N__24676\
        );

    \I__2801\ : Odrv12
    port map (
            O => \N__24676\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\
        );

    \I__2800\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24670\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__24670\,
            I => \phase_controller_inst2.stoper_tr.counter_i_14\
        );

    \I__2798\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24664\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__24664\,
            I => \N__24661\
        );

    \I__2796\ : Odrv12
    port map (
            O => \N__24661\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__24658\,
            I => \N__24655\
        );

    \I__2794\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24652\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__24652\,
            I => \phase_controller_inst2.stoper_tr.counter_i_15\
        );

    \I__2792\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24646\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24643\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__24643\,
            I => \N__24640\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__24640\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt16\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__24637\,
            I => \N__24634\
        );

    \I__2787\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24631\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24628\
        );

    \I__2785\ : Span4Mux_h
    port map (
            O => \N__24628\,
            I => \N__24625\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__24625\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\
        );

    \I__2783\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24619\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__24619\,
            I => \N__24616\
        );

    \I__2781\ : Span4Mux_h
    port map (
            O => \N__24616\,
            I => \N__24613\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__24613\,
            I => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__24610\,
            I => \N__24607\
        );

    \I__2778\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24604\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__24601\,
            I => \N__24598\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__24598\,
            I => \phase_controller_inst2.stoper_tr.un6_running_lt18\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__24595\,
            I => \N__24592\
        );

    \I__2773\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24589\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__24586\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\
        );

    \I__2770\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__24580\,
            I => \phase_controller_inst2.stoper_tr.counter_i_2\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__24577\,
            I => \N__24574\
        );

    \I__2767\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24571\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24568\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__24568\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\
        );

    \I__2764\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__24562\,
            I => \phase_controller_inst2.stoper_tr.counter_i_3\
        );

    \I__2762\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24556\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__24556\,
            I => \N__24553\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__24553\,
            I => \N__24550\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__24547\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__2756\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24538\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__24538\,
            I => \phase_controller_inst2.stoper_tr.counter_i_4\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__24535\,
            I => \N__24532\
        );

    \I__2753\ : InMux
    port map (
            O => \N__24532\,
            I => \N__24529\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__24529\,
            I => \N__24526\
        );

    \I__2751\ : Odrv12
    port map (
            O => \N__24526\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\
        );

    \I__2750\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24520\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__24520\,
            I => \phase_controller_inst2.stoper_tr.counter_i_5\
        );

    \I__2748\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__24514\,
            I => \N__24511\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__24511\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__2744\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24502\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__24502\,
            I => \phase_controller_inst2.stoper_tr.counter_i_6\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__24499\,
            I => \N__24496\
        );

    \I__2741\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24493\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24490\
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__24490\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\
        );

    \I__2738\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__24484\,
            I => \phase_controller_inst2.stoper_tr.counter_i_7\
        );

    \I__2736\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__24475\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__24472\,
            I => \N__24469\
        );

    \I__2732\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24466\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__24466\,
            I => \phase_controller_inst2.stoper_tr.counter_i_8\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__24463\,
            I => \N__24460\
        );

    \I__2729\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24457\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__24457\,
            I => \N__24454\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__24454\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\
        );

    \I__2726\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24448\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__24448\,
            I => \phase_controller_inst2.stoper_tr.counter_i_9\
        );

    \I__2724\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24439\
        );

    \I__2723\ : InMux
    port map (
            O => \N__24444\,
            I => \N__24439\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__24439\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\
        );

    \I__2721\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24430\
        );

    \I__2720\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24430\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__24430\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\
        );

    \I__2718\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24421\
        );

    \I__2717\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24421\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__24421\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\
        );

    \I__2715\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24412\
        );

    \I__2714\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24412\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__24412\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\
        );

    \I__2712\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24406\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__24406\,
            I => \N__24403\
        );

    \I__2710\ : Odrv12
    port map (
            O => \N__24403\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__24400\,
            I => \N__24397\
        );

    \I__2708\ : InMux
    port map (
            O => \N__24397\,
            I => \N__24394\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__24394\,
            I => \phase_controller_inst2.stoper_tr.counter_i_0\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__24391\,
            I => \N__24388\
        );

    \I__2705\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__2703\ : Odrv12
    port map (
            O => \N__24382\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\
        );

    \I__2702\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__24376\,
            I => \phase_controller_inst2.stoper_tr.counter_i_1\
        );

    \I__2700\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24343\
        );

    \I__2699\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24343\
        );

    \I__2698\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24343\
        );

    \I__2697\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24343\
        );

    \I__2696\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24330\
        );

    \I__2695\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24330\
        );

    \I__2694\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24321\
        );

    \I__2693\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24321\
        );

    \I__2692\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24321\
        );

    \I__2691\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24321\
        );

    \I__2690\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24312\
        );

    \I__2689\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24312\
        );

    \I__2688\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24312\
        );

    \I__2687\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24312\
        );

    \I__2686\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24303\
        );

    \I__2685\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24303\
        );

    \I__2684\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24303\
        );

    \I__2683\ : InMux
    port map (
            O => \N__24356\,
            I => \N__24303\
        );

    \I__2682\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24294\
        );

    \I__2681\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24294\
        );

    \I__2680\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24294\
        );

    \I__2679\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24294\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__24343\,
            I => \N__24291\
        );

    \I__2677\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24282\
        );

    \I__2676\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24282\
        );

    \I__2675\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24282\
        );

    \I__2674\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24282\
        );

    \I__2673\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24273\
        );

    \I__2672\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24273\
        );

    \I__2671\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24273\
        );

    \I__2670\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24273\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__24330\,
            I => \N__24268\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24268\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__24312\,
            I => \N__24257\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__24303\,
            I => \N__24257\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24257\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__24291\,
            I => \N__24257\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24257\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24254\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__24268\,
            I => \N__24249\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__24257\,
            I => \N__24249\
        );

    \I__2659\ : Odrv12
    port map (
            O => \N__24254\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__24249\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__2657\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24241\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__24241\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__24238\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\
        );

    \I__2654\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24232\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__24232\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__24229\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\
        );

    \I__2651\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24223\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__24223\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__24220\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\
        );

    \I__2648\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24213\
        );

    \I__2647\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24210\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__24213\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__24210\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__2644\ : InMux
    port map (
            O => \N__24205\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__2643\ : InMux
    port map (
            O => \N__24202\,
            I => \bfn_7_10_0_\
        );

    \I__2642\ : InMux
    port map (
            O => \N__24199\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__2641\ : InMux
    port map (
            O => \N__24196\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__2640\ : InMux
    port map (
            O => \N__24193\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__2639\ : InMux
    port map (
            O => \N__24190\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__2638\ : InMux
    port map (
            O => \N__24187\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__2637\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24181\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__24181\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__24178\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__2634\ : InMux
    port map (
            O => \N__24175\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__2633\ : InMux
    port map (
            O => \N__24172\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__2632\ : InMux
    port map (
            O => \N__24169\,
            I => \bfn_7_9_0_\
        );

    \I__2631\ : InMux
    port map (
            O => \N__24166\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__2630\ : InMux
    port map (
            O => \N__24163\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__2629\ : InMux
    port map (
            O => \N__24160\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__2628\ : InMux
    port map (
            O => \N__24157\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__2627\ : InMux
    port map (
            O => \N__24154\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__2626\ : InMux
    port map (
            O => \N__24151\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__2625\ : InMux
    port map (
            O => \N__24148\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__2624\ : InMux
    port map (
            O => \N__24145\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__2623\ : InMux
    port map (
            O => \N__24142\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__2622\ : InMux
    port map (
            O => \N__24139\,
            I => \bfn_7_8_0_\
        );

    \I__2621\ : InMux
    port map (
            O => \N__24136\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__2620\ : InMux
    port map (
            O => \N__24133\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__2619\ : InMux
    port map (
            O => \N__24130\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__2618\ : InMux
    port map (
            O => \N__24127\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__2617\ : InMux
    port map (
            O => \N__24124\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__2616\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24115\
        );

    \I__2615\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24115\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24112\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__24112\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\
        );

    \I__2612\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24103\
        );

    \I__2611\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24103\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__24100\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\
        );

    \I__2608\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24091\
        );

    \I__2607\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24091\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24088\
        );

    \I__2605\ : Odrv12
    port map (
            O => \N__24088\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\
        );

    \I__2604\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24079\
        );

    \I__2603\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24079\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__24079\,
            I => \N__24076\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__24076\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\
        );

    \I__2600\ : InMux
    port map (
            O => \N__24073\,
            I => \bfn_7_7_0_\
        );

    \I__2599\ : InMux
    port map (
            O => \N__24070\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__2598\ : InMux
    port map (
            O => \N__24067\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__2597\ : InMux
    port map (
            O => \N__24064\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__2596\ : InMux
    port map (
            O => \N__24061\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__2595\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24052\
        );

    \I__2594\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24052\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__24052\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\
        );

    \I__2592\ : InMux
    port map (
            O => \N__24049\,
            I => \N__24043\
        );

    \I__2591\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24043\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__24043\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__24040\,
            I => \N__24036\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__24039\,
            I => \N__24033\
        );

    \I__2587\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24028\
        );

    \I__2586\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24028\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__24028\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\
        );

    \I__2584\ : InMux
    port map (
            O => \N__24025\,
            I => \N__24019\
        );

    \I__2583\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24019\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__24019\,
            I => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\
        );

    \I__2581\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24010\
        );

    \I__2580\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24010\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__24010\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\
        );

    \I__2578\ : InMux
    port map (
            O => \N__24007\,
            I => \N__24001\
        );

    \I__2577\ : InMux
    port map (
            O => \N__24006\,
            I => \N__24001\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__24001\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__23998\,
            I => \N__23994\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__23997\,
            I => \N__23991\
        );

    \I__2573\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23986\
        );

    \I__2572\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23986\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__23986\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\
        );

    \I__2570\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23977\
        );

    \I__2569\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23977\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__23977\,
            I => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\
        );

    \I__2567\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23969\
        );

    \I__2566\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23966\
        );

    \I__2565\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23963\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__23969\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__23966\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__23963\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__2561\ : InMux
    port map (
            O => \N__23956\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__2560\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23948\
        );

    \I__2559\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23945\
        );

    \I__2558\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23942\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__23948\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__23945\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__23942\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__2554\ : InMux
    port map (
            O => \N__23935\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__2553\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23927\
        );

    \I__2552\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23924\
        );

    \I__2551\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23921\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__23927\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__23924\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__23921\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__2547\ : InMux
    port map (
            O => \N__23914\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__2546\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23906\
        );

    \I__2545\ : InMux
    port map (
            O => \N__23910\,
            I => \N__23903\
        );

    \I__2544\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23900\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__23906\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__23903\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__23900\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__2540\ : InMux
    port map (
            O => \N__23893\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__2539\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23885\
        );

    \I__2538\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23882\
        );

    \I__2537\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23879\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__23885\,
            I => \N__23876\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__23882\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__23879\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__23876\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__2532\ : InMux
    port map (
            O => \N__23869\,
            I => \bfn_4_19_0_\
        );

    \I__2531\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23852\
        );

    \I__2530\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23852\
        );

    \I__2529\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23843\
        );

    \I__2528\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23843\
        );

    \I__2527\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23843\
        );

    \I__2526\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23843\
        );

    \I__2525\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23834\
        );

    \I__2524\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23834\
        );

    \I__2523\ : InMux
    port map (
            O => \N__23858\,
            I => \N__23834\
        );

    \I__2522\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23834\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23831\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__23843\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__23834\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__23831\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__2517\ : InMux
    port map (
            O => \N__23824\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__2516\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23816\
        );

    \I__2515\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23813\
        );

    \I__2514\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23810\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23807\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__23813\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__23810\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__23807\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__2509\ : InMux
    port map (
            O => \N__23800\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2508\ : IoInMux
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__23794\,
            I => \N__23791\
        );

    \I__2506\ : Span4Mux_s3_v
    port map (
            O => \N__23791\,
            I => \N__23788\
        );

    \I__2505\ : Sp12to4
    port map (
            O => \N__23788\,
            I => \N__23785\
        );

    \I__2504\ : Span12Mux_s10_h
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__2503\ : Span12Mux_h
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__2502\ : Span12Mux_v
    port map (
            O => \N__23779\,
            I => \N__23776\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__23776\,
            I => pwm_output_c
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__23773\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2499\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23767\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__23767\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__23764\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__2496\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23756\
        );

    \I__2495\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23753\
        );

    \I__2494\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23750\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__23756\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__23753\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__23750\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__2490\ : InMux
    port map (
            O => \N__23743\,
            I => \bfn_4_18_0_\
        );

    \I__2489\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23735\
        );

    \I__2488\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23732\
        );

    \I__2487\ : InMux
    port map (
            O => \N__23738\,
            I => \N__23729\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__23735\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__23732\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__23729\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__2483\ : InMux
    port map (
            O => \N__23722\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__2482\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23714\
        );

    \I__2481\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23711\
        );

    \I__2480\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23708\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__23714\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__23711\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__23708\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__2476\ : InMux
    port map (
            O => \N__23701\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__2475\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23693\
        );

    \I__2474\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23690\
        );

    \I__2473\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23687\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__23693\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__23690\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__23687\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__2469\ : InMux
    port map (
            O => \N__23680\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__23677\,
            I => \N__23674\
        );

    \I__2467\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23671\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__23665\,
            I => \pwm_generator_inst.N_181_i\
        );

    \I__2463\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23659\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__23659\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__23656\,
            I => \N__23653\
        );

    \I__2460\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23647\
        );

    \I__2458\ : Span12Mux_h
    port map (
            O => \N__23647\,
            I => \N__23644\
        );

    \I__2457\ : Odrv12
    port map (
            O => \N__23644\,
            I => \pwm_generator_inst.N_182_i\
        );

    \I__2456\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23638\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__23638\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__23635\,
            I => \N__23632\
        );

    \I__2453\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23629\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__23626\,
            I => \N__23623\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__23623\,
            I => \pwm_generator_inst.N_183_i\
        );

    \I__2449\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23617\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__23617\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2447\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23611\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__23611\,
            I => \pwm_generator_inst.N_184_i\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__23608\,
            I => \N__23605\
        );

    \I__2444\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23602\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__23602\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__23599\,
            I => \N__23596\
        );

    \I__2441\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23593\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__23593\,
            I => \N__23590\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__23590\,
            I => \N__23587\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__23587\,
            I => \pwm_generator_inst.N_185_i\
        );

    \I__2437\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23581\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__23581\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__23578\,
            I => \N__23575\
        );

    \I__2434\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23572\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__23572\,
            I => \N__23569\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__23569\,
            I => \pwm_generator_inst.N_186_i\
        );

    \I__2431\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23563\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__23563\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__23560\,
            I => \N__23557\
        );

    \I__2428\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23554\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__23554\,
            I => \pwm_generator_inst.N_187_i\
        );

    \I__2426\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23548\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__23548\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23542\
        );

    \I__2423\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23539\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__23536\,
            I => \N__23533\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__23533\,
            I => \pwm_generator_inst.N_188_i\
        );

    \I__2419\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23527\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__23527\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__23524\,
            I => \N__23520\
        );

    \I__2416\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23517\
        );

    \I__2415\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23514\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__23517\,
            I => \pwm_generator_inst.un18_threshold1_24\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__23514\,
            I => \pwm_generator_inst.un18_threshold1_24\
        );

    \I__2412\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23506\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__23506\,
            I => \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO\
        );

    \I__2410\ : InMux
    port map (
            O => \N__23503\,
            I => \pwm_generator_inst.un22_threshold_1_cry_6\
        );

    \I__2409\ : InMux
    port map (
            O => \N__23500\,
            I => \bfn_2_18_0_\
        );

    \I__2408\ : InMux
    port map (
            O => \N__23497\,
            I => \pwm_generator_inst.un22_threshold_1_cry_8\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__2406\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23488\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__23488\,
            I => \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO\
        );

    \I__2404\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23482\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23478\
        );

    \I__2402\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23475\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__23478\,
            I => \pwm_generator_inst.un22_threshold_1\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__23475\,
            I => \pwm_generator_inst.un22_threshold_1\
        );

    \I__2399\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23466\
        );

    \I__2398\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23463\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__23466\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__23463\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\
        );

    \I__2395\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23454\
        );

    \I__2394\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23451\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23448\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23445\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__23448\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__23445\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__23440\,
            I => \N__23436\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__23439\,
            I => \N__23433\
        );

    \I__2387\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23428\
        );

    \I__2386\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23428\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__23428\,
            I => \pwm_generator_inst.un18_threshold1_25\
        );

    \I__2384\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23422\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__23422\,
            I => \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO\
        );

    \I__2382\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__23416\,
            I => \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO\
        );

    \I__2380\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23409\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__23412\,
            I => \N__23406\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23403\
        );

    \I__2377\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23400\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__23403\,
            I => \pwm_generator_inst.un18_threshold1_18\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__23400\,
            I => \pwm_generator_inst.un18_threshold1_18\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__23395\,
            I => \N__23388\
        );

    \I__2373\ : InMux
    port map (
            O => \N__23394\,
            I => \N__23380\
        );

    \I__2372\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23375\
        );

    \I__2371\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23375\
        );

    \I__2370\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23368\
        );

    \I__2369\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23368\
        );

    \I__2368\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23368\
        );

    \I__2367\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23359\
        );

    \I__2366\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23359\
        );

    \I__2365\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23359\
        );

    \I__2364\ : InMux
    port map (
            O => \N__23383\,
            I => \N__23359\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23350\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__23375\,
            I => \N__23350\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N__23350\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__23359\,
            I => \N__23350\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__23350\,
            I => \N__23347\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__23347\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\
        );

    \I__2357\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23340\
        );

    \I__2356\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23337\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__23340\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__23337\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__23332\,
            I => \N__23329\
        );

    \I__2352\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23326\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__23326\,
            I => \pwm_generator_inst.N_179_i\
        );

    \I__2350\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23320\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__23320\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__23317\,
            I => \N__23314\
        );

    \I__2347\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23311\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__23311\,
            I => \pwm_generator_inst.N_180_i\
        );

    \I__2345\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23305\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__23305\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__23302\,
            I => \N__23299\
        );

    \I__2342\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23296\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__23296\,
            I => \N__23292\
        );

    \I__2340\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23289\
        );

    \I__2339\ : Span4Mux_h
    port map (
            O => \N__23292\,
            I => \N__23284\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23284\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__23284\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\
        );

    \I__2336\ : InMux
    port map (
            O => \N__23281\,
            I => \pwm_generator_inst.un22_threshold_1_cry_0\
        );

    \I__2335\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23274\
        );

    \I__2334\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23271\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__23274\,
            I => \pwm_generator_inst.un18_threshold1_19\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__23271\,
            I => \pwm_generator_inst.un18_threshold1_19\
        );

    \I__2331\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23263\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__23263\,
            I => \N__23260\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__23260\,
            I => \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO\
        );

    \I__2328\ : InMux
    port map (
            O => \N__23257\,
            I => \pwm_generator_inst.un22_threshold_1_cry_1\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__23254\,
            I => \N__23250\
        );

    \I__2326\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23247\
        );

    \I__2325\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23244\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__23247\,
            I => \pwm_generator_inst.un18_threshold1_20\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__23244\,
            I => \pwm_generator_inst.un18_threshold1_20\
        );

    \I__2322\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23236\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__23233\,
            I => \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO\
        );

    \I__2319\ : InMux
    port map (
            O => \N__23230\,
            I => \pwm_generator_inst.un22_threshold_1_cry_2\
        );

    \I__2318\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23223\
        );

    \I__2317\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23220\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__23223\,
            I => \pwm_generator_inst.un18_threshold1_21\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__23220\,
            I => \pwm_generator_inst.un18_threshold1_21\
        );

    \I__2314\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23209\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__23209\,
            I => \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO\
        );

    \I__2311\ : InMux
    port map (
            O => \N__23206\,
            I => \pwm_generator_inst.un22_threshold_1_cry_3\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__23203\,
            I => \N__23199\
        );

    \I__2309\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23196\
        );

    \I__2308\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23193\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__23196\,
            I => \pwm_generator_inst.un18_threshold1_22\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__23193\,
            I => \pwm_generator_inst.un18_threshold1_22\
        );

    \I__2305\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__23185\,
            I => \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO\
        );

    \I__2303\ : InMux
    port map (
            O => \N__23182\,
            I => \pwm_generator_inst.un22_threshold_1_cry_4\
        );

    \I__2302\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23175\
        );

    \I__2301\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23172\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__23175\,
            I => \pwm_generator_inst.un18_threshold1_23\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__23172\,
            I => \pwm_generator_inst.un18_threshold1_23\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__23167\,
            I => \N__23164\
        );

    \I__2297\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23161\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__23161\,
            I => \N__23158\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__23158\,
            I => \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO\
        );

    \I__2294\ : InMux
    port map (
            O => \N__23155\,
            I => \pwm_generator_inst.un22_threshold_1_cry_5\
        );

    \I__2293\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__23149\,
            I => \N__23146\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__23146\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7\
        );

    \I__2290\ : InMux
    port map (
            O => \N__23143\,
            I => \bfn_1_25_0_\
        );

    \I__2289\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__23137\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7\
        );

    \I__2287\ : InMux
    port map (
            O => \N__23134\,
            I => \pwm_generator_inst.un3_threshold_cry_16\
        );

    \I__2286\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23128\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__23128\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0\
        );

    \I__2284\ : InMux
    port map (
            O => \N__23125\,
            I => \pwm_generator_inst.un3_threshold_cry_17\
        );

    \I__2283\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23118\
        );

    \I__2282\ : InMux
    port map (
            O => \N__23121\,
            I => \N__23115\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__23118\,
            I => \N__23110\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__23115\,
            I => \N__23110\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__23110\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\
        );

    \I__2278\ : InMux
    port map (
            O => \N__23107\,
            I => \pwm_generator_inst.un3_threshold_cry_18\
        );

    \I__2277\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__23092\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__2272\ : InMux
    port map (
            O => \N__23089\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__2271\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23083\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__23083\,
            I => \N__23080\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__23080\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__2267\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__23071\,
            I => \N__23067\
        );

    \I__2265\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23064\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__23067\,
            I => \N__23059\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23059\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__23059\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__2260\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23050\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__23050\,
            I => \N__23047\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__23047\,
            I => \N__23043\
        );

    \I__2257\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23040\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__23043\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__23040\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__2253\ : InMux
    port map (
            O => \N__23032\,
            I => \N__23029\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__23029\,
            I => \N__23025\
        );

    \I__2251\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23022\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__23025\,
            I => \N__23019\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__23022\,
            I => \N__23016\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__23019\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__23016\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\
        );

    \I__2246\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23008\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__23004\
        );

    \I__2244\ : InMux
    port map (
            O => \N__23007\,
            I => \N__23001\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__23004\,
            I => \N__22998\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22995\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__22998\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__22995\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\
        );

    \I__2239\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__22987\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0\
        );

    \I__2237\ : InMux
    port map (
            O => \N__22984\,
            I => \bfn_1_24_0_\
        );

    \I__2236\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__22978\,
            I => \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8\
        );

    \I__2234\ : InMux
    port map (
            O => \N__22975\,
            I => \pwm_generator_inst.un3_threshold_cry_8\
        );

    \I__2233\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22969\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__22969\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8\
        );

    \I__2231\ : InMux
    port map (
            O => \N__22966\,
            I => \pwm_generator_inst.un3_threshold_cry_9\
        );

    \I__2230\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22960\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__22960\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7\
        );

    \I__2228\ : InMux
    port map (
            O => \N__22957\,
            I => \pwm_generator_inst.un3_threshold_cry_10\
        );

    \I__2227\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__22951\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7\
        );

    \I__2225\ : InMux
    port map (
            O => \N__22948\,
            I => \pwm_generator_inst.un3_threshold_cry_11\
        );

    \I__2224\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22942\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__22942\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7\
        );

    \I__2222\ : InMux
    port map (
            O => \N__22939\,
            I => \pwm_generator_inst.un3_threshold_cry_12\
        );

    \I__2221\ : InMux
    port map (
            O => \N__22936\,
            I => \N__22933\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__22933\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7\
        );

    \I__2219\ : InMux
    port map (
            O => \N__22930\,
            I => \pwm_generator_inst.un3_threshold_cry_13\
        );

    \I__2218\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22924\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__22924\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7\
        );

    \I__2216\ : InMux
    port map (
            O => \N__22921\,
            I => \pwm_generator_inst.un3_threshold_cry_14\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__2214\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22912\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__22912\,
            I => \N__22909\
        );

    \I__2212\ : Span12Mux_v
    port map (
            O => \N__22909\,
            I => \N__22906\
        );

    \I__2211\ : Span12Mux_h
    port map (
            O => \N__22906\,
            I => \N__22903\
        );

    \I__2210\ : Span12Mux_h
    port map (
            O => \N__22903\,
            I => \N__22900\
        );

    \I__2209\ : Odrv12
    port map (
            O => \N__22900\,
            I => \pwm_generator_inst.O_0_8\
        );

    \I__2208\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__2206\ : Span12Mux_s1_h
    port map (
            O => \N__22891\,
            I => \N__22888\
        );

    \I__2205\ : Odrv12
    port map (
            O => \N__22888\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0\
        );

    \I__2204\ : InMux
    port map (
            O => \N__22885\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__2202\ : InMux
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__22876\,
            I => \N__22873\
        );

    \I__2200\ : Span12Mux_v
    port map (
            O => \N__22873\,
            I => \N__22870\
        );

    \I__2199\ : Span12Mux_h
    port map (
            O => \N__22870\,
            I => \N__22867\
        );

    \I__2198\ : Span12Mux_h
    port map (
            O => \N__22867\,
            I => \N__22864\
        );

    \I__2197\ : Odrv12
    port map (
            O => \N__22864\,
            I => \pwm_generator_inst.O_0_9\
        );

    \I__2196\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22858\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__22858\,
            I => \N__22855\
        );

    \I__2194\ : Sp12to4
    port map (
            O => \N__22855\,
            I => \N__22852\
        );

    \I__2193\ : Odrv12
    port map (
            O => \N__22852\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0\
        );

    \I__2192\ : InMux
    port map (
            O => \N__22849\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__2191\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__22843\,
            I => \N__22840\
        );

    \I__2189\ : Span4Mux_v
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__22837\,
            I => \N__22834\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__22834\,
            I => \N__22831\
        );

    \I__2186\ : Sp12to4
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__2185\ : Span12Mux_h
    port map (
            O => \N__22828\,
            I => \N__22825\
        );

    \I__2184\ : Odrv12
    port map (
            O => \N__22825\,
            I => \pwm_generator_inst.O_0_10\
        );

    \I__2183\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22819\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__22819\,
            I => \N__22816\
        );

    \I__2181\ : Span4Mux_v
    port map (
            O => \N__22816\,
            I => \N__22813\
        );

    \I__2180\ : Span4Mux_v
    port map (
            O => \N__22813\,
            I => \N__22810\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__22810\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0\
        );

    \I__2178\ : InMux
    port map (
            O => \N__22807\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__2177\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22801\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__22801\,
            I => \N__22798\
        );

    \I__2175\ : Span12Mux_s11_v
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__2174\ : Span12Mux_h
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__2173\ : Span12Mux_h
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__22789\,
            I => \pwm_generator_inst.O_0_11\
        );

    \I__2171\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22783\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__22780\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0\
        );

    \I__2168\ : InMux
    port map (
            O => \N__22777\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__2167\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__22771\,
            I => \N__22768\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__22765\,
            I => \N__22762\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__2162\ : Sp12to4
    port map (
            O => \N__22759\,
            I => \N__22756\
        );

    \I__2161\ : Span12Mux_h
    port map (
            O => \N__22756\,
            I => \N__22753\
        );

    \I__2160\ : Odrv12
    port map (
            O => \N__22753\,
            I => \pwm_generator_inst.O_0_12\
        );

    \I__2159\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__2157\ : Span4Mux_s1_h
    port map (
            O => \N__22744\,
            I => \N__22741\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__22741\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0\
        );

    \I__2155\ : InMux
    port map (
            O => \N__22738\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__2154\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22732\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22729\
        );

    \I__2152\ : Span12Mux_s9_v
    port map (
            O => \N__22729\,
            I => \N__22726\
        );

    \I__2151\ : Span12Mux_h
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__2150\ : Span12Mux_h
    port map (
            O => \N__22723\,
            I => \N__22720\
        );

    \I__2149\ : Odrv12
    port map (
            O => \N__22720\,
            I => \pwm_generator_inst.O_0_13\
        );

    \I__2148\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22714\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22711\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__22711\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0\
        );

    \I__2145\ : InMux
    port map (
            O => \N__22708\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__2144\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22702\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22699\
        );

    \I__2142\ : Span12Mux_s8_v
    port map (
            O => \N__22699\,
            I => \N__22696\
        );

    \I__2141\ : Span12Mux_h
    port map (
            O => \N__22696\,
            I => \N__22693\
        );

    \I__2140\ : Span12Mux_h
    port map (
            O => \N__22693\,
            I => \N__22690\
        );

    \I__2139\ : Odrv12
    port map (
            O => \N__22690\,
            I => \pwm_generator_inst.O_0_14\
        );

    \I__2138\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22684\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__22684\,
            I => \N__22681\
        );

    \I__2136\ : Span4Mux_s1_h
    port map (
            O => \N__22681\,
            I => \N__22678\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__22678\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0\
        );

    \I__2134\ : InMux
    port map (
            O => \N__22675\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__22672\,
            I => \N__22669\
        );

    \I__2132\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22666\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__22666\,
            I => \N__22663\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__22663\,
            I => \N__22660\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__22660\,
            I => \pwm_generator_inst.un5_threshold_2_11\
        );

    \I__2128\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__22651\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0\
        );

    \I__2125\ : InMux
    port map (
            O => \N__22648\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_10\
        );

    \I__2124\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22642\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__22642\,
            I => \N__22639\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__22636\,
            I => \pwm_generator_inst.un5_threshold_2_12\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__22633\,
            I => \N__22630\
        );

    \I__2119\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22627\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22624\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__22624\,
            I => \N__22621\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__22621\,
            I => \pwm_generator_inst.un5_threshold_2_13\
        );

    \I__2115\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22615\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22612\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__22612\,
            I => \N__22609\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__22609\,
            I => \pwm_generator_inst.un5_threshold_2_14\
        );

    \I__2111\ : InMux
    port map (
            O => \N__22606\,
            I => \bfn_1_21_0_\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__2109\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__22594\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__22591\,
            I => \N__22584\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__22590\,
            I => \N__22580\
        );

    \I__2104\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22576\
        );

    \I__2103\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22573\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22562\
        );

    \I__2101\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22562\
        );

    \I__2100\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22562\
        );

    \I__2099\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22562\
        );

    \I__2098\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22562\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__22576\,
            I => \N__22557\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__22573\,
            I => \N__22557\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22552\
        );

    \I__2094\ : Span4Mux_v
    port map (
            O => \N__22557\,
            I => \N__22552\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__22552\,
            I => \N__22549\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__22549\,
            I => \pwm_generator_inst.un5_threshold_1_26\
        );

    \I__2091\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22543\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__22540\,
            I => \pwm_generator_inst.un5_threshold_2_1_16\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__22537\,
            I => \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22530\
        );

    \I__2086\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22527\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__22530\,
            I => \N__22524\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__22527\,
            I => \N__22521\
        );

    \I__2083\ : Span4Mux_h
    port map (
            O => \N__22524\,
            I => \N__22518\
        );

    \I__2082\ : Span4Mux_h
    port map (
            O => \N__22521\,
            I => \N__22515\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__22518\,
            I => \pwm_generator_inst.un5_threshold_2_1_15\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__22515\,
            I => \pwm_generator_inst.un5_threshold_2_1_15\
        );

    \I__2079\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__22507\,
            I => \pwm_generator_inst.un5_threshold_add_1_axb_16\
        );

    \I__2077\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__22498\,
            I => \N__22495\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__22495\,
            I => \pwm_generator_inst.un5_threshold_1_19\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__22492\,
            I => \N__22489\
        );

    \I__2072\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22486\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22483\
        );

    \I__2070\ : Span4Mux_h
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__22480\,
            I => \pwm_generator_inst.un5_threshold_2_4\
        );

    \I__2068\ : InMux
    port map (
            O => \N__22477\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_3\
        );

    \I__2067\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__22468\,
            I => \N__22465\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__22465\,
            I => \pwm_generator_inst.un5_threshold_1_20\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__22462\,
            I => \N__22459\
        );

    \I__2062\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__22453\,
            I => \N__22450\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__22450\,
            I => \pwm_generator_inst.un5_threshold_2_5\
        );

    \I__2058\ : InMux
    port map (
            O => \N__22447\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_4\
        );

    \I__2057\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22441\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__22438\,
            I => \N__22435\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__22435\,
            I => \pwm_generator_inst.un5_threshold_1_21\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__2052\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22426\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__22420\,
            I => \pwm_generator_inst.un5_threshold_2_6\
        );

    \I__2048\ : InMux
    port map (
            O => \N__22417\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_5\
        );

    \I__2047\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__22405\,
            I => \pwm_generator_inst.un5_threshold_1_22\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \N__22399\
        );

    \I__2042\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22396\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22393\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__22390\,
            I => \pwm_generator_inst.un5_threshold_2_7\
        );

    \I__2038\ : InMux
    port map (
            O => \N__22387\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_6\
        );

    \I__2037\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22381\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__22381\,
            I => \N__22378\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__22378\,
            I => \N__22375\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__22375\,
            I => \N__22372\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__22372\,
            I => \pwm_generator_inst.un5_threshold_1_23\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__22369\,
            I => \N__22366\
        );

    \I__2031\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22363\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__22363\,
            I => \N__22360\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__22357\,
            I => \pwm_generator_inst.un5_threshold_2_8\
        );

    \I__2027\ : InMux
    port map (
            O => \N__22354\,
            I => \bfn_1_20_0_\
        );

    \I__2026\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22348\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__22339\,
            I => \pwm_generator_inst.un5_threshold_1_24\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__22336\,
            I => \N__22333\
        );

    \I__2020\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22330\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__2018\ : Span4Mux_h
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__22324\,
            I => \pwm_generator_inst.un5_threshold_2_9\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__2015\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22314\
        );

    \I__2014\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22311\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__22314\,
            I => \N__22308\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22305\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__22308\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__22305\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\
        );

    \I__2009\ : InMux
    port map (
            O => \N__22300\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_8\
        );

    \I__2008\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22294\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__22291\,
            I => \N__22288\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__22285\,
            I => \pwm_generator_inst.un5_threshold_1_25\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__2002\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22276\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__22273\,
            I => \N__22270\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__22270\,
            I => \pwm_generator_inst.un5_threshold_2_10\
        );

    \I__1998\ : InMux
    port map (
            O => \N__22267\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_9\
        );

    \I__1997\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22261\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22258\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__22258\,
            I => \pwm_generator_inst.un18_threshold_1_axb_17\
        );

    \I__1994\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22252\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__22252\,
            I => \pwm_generator_inst.un18_threshold_1_axb_25\
        );

    \I__1992\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22246\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__22246\,
            I => \N__22243\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__22243\,
            I => \pwm_generator_inst.un18_threshold_1_axb_20\
        );

    \I__1989\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__22237\,
            I => \pwm_generator_inst.un18_threshold_1_axb_24\
        );

    \I__1987\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22231\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__22228\,
            I => \pwm_generator_inst.un18_threshold_1_axb_18\
        );

    \I__1984\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22222\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__22222\,
            I => \N__22219\
        );

    \I__1982\ : Span4Mux_h
    port map (
            O => \N__22219\,
            I => \N__22216\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__22216\,
            I => \pwm_generator_inst.un5_threshold_2_0\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__22213\,
            I => \N__22210\
        );

    \I__1979\ : InMux
    port map (
            O => \N__22210\,
            I => \N__22207\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22204\
        );

    \I__1977\ : Span12Mux_v
    port map (
            O => \N__22204\,
            I => \N__22201\
        );

    \I__1976\ : Odrv12
    port map (
            O => \N__22201\,
            I => \pwm_generator_inst.un5_threshold_1_15\
        );

    \I__1975\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22195\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__22195\,
            I => \N__22192\
        );

    \I__1973\ : Odrv12
    port map (
            O => \N__22192\,
            I => \pwm_generator_inst.un18_threshold_1_axb_15\
        );

    \I__1972\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__22186\,
            I => \N__22183\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__22183\,
            I => \N__22180\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__22180\,
            I => \pwm_generator_inst.un5_threshold_2_1\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__22177\,
            I => \N__22174\
        );

    \I__1967\ : InMux
    port map (
            O => \N__22174\,
            I => \N__22171\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__22168\,
            I => \N__22165\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__22162\,
            I => \pwm_generator_inst.un5_threshold_1_16\
        );

    \I__1962\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22156\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__22156\,
            I => \N__22153\
        );

    \I__1960\ : Odrv12
    port map (
            O => \N__22153\,
            I => \pwm_generator_inst.un18_threshold_1_axb_16\
        );

    \I__1959\ : InMux
    port map (
            O => \N__22150\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_0\
        );

    \I__1958\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22144\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__22141\,
            I => \N__22138\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__22138\,
            I => \pwm_generator_inst.un5_threshold_2_2\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__1953\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__22126\,
            I => \N__22123\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__22120\,
            I => \pwm_generator_inst.un5_threshold_1_17\
        );

    \I__1948\ : InMux
    port map (
            O => \N__22117\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_1\
        );

    \I__1947\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22108\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__22108\,
            I => \N__22105\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__22105\,
            I => \pwm_generator_inst.un5_threshold_2_3\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__1942\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__22093\,
            I => \N__22090\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__22090\,
            I => \pwm_generator_inst.un5_threshold_1_18\
        );

    \I__1938\ : InMux
    port map (
            O => \N__22087\,
            I => \pwm_generator_inst.un5_threshold_add_1_cry_2\
        );

    \I__1937\ : InMux
    port map (
            O => \N__22084\,
            I => \pwm_generator_inst.un18_threshold_1_cry_22\
        );

    \I__1936\ : InMux
    port map (
            O => \N__22081\,
            I => \bfn_1_17_0_\
        );

    \I__1935\ : InMux
    port map (
            O => \N__22078\,
            I => \pwm_generator_inst.un18_threshold_1_cry_24\
        );

    \I__1934\ : InMux
    port map (
            O => \N__22075\,
            I => \pwm_generator_inst.un18_threshold_1_cry_25\
        );

    \I__1933\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22069\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__22069\,
            I => \pwm_generator_inst.un18_threshold_1_axb_19\
        );

    \I__1931\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22063\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__22063\,
            I => \pwm_generator_inst.un18_threshold_1_axb_21\
        );

    \I__1929\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__22057\,
            I => \pwm_generator_inst.un18_threshold_1_axb_22\
        );

    \I__1927\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22051\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__22051\,
            I => \pwm_generator_inst.un18_threshold_1_axb_23\
        );

    \I__1925\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__22045\,
            I => \N__22042\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__22042\,
            I => \N__22039\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__22039\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1921\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22033\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__22033\,
            I => \pwm_generator_inst.un18_threshold_1_axb_14\
        );

    \I__1919\ : InMux
    port map (
            O => \N__22030\,
            I => \pwm_generator_inst.un18_threshold_1_cry_16\
        );

    \I__1918\ : InMux
    port map (
            O => \N__22027\,
            I => \pwm_generator_inst.un18_threshold_1_cry_17\
        );

    \I__1917\ : InMux
    port map (
            O => \N__22024\,
            I => \pwm_generator_inst.un18_threshold_1_cry_18\
        );

    \I__1916\ : InMux
    port map (
            O => \N__22021\,
            I => \pwm_generator_inst.un18_threshold_1_cry_19\
        );

    \I__1915\ : InMux
    port map (
            O => \N__22018\,
            I => \pwm_generator_inst.un18_threshold_1_cry_20\
        );

    \I__1914\ : InMux
    port map (
            O => \N__22015\,
            I => \pwm_generator_inst.un18_threshold_1_cry_21\
        );

    \I__1913\ : InMux
    port map (
            O => \N__22012\,
            I => \N__22009\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__22003\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1909\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__21997\,
            I => \pwm_generator_inst.un18_threshold_1_axb_6\
        );

    \I__1907\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21991\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21988\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__21988\,
            I => \N__21985\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__21985\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1903\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21979\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__21979\,
            I => \pwm_generator_inst.un18_threshold_1_axb_7\
        );

    \I__1901\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21973\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__21973\,
            I => \N__21970\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__21970\,
            I => \N__21967\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__21967\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1897\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__21961\,
            I => \pwm_generator_inst.un18_threshold_1_axb_8\
        );

    \I__1895\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21955\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__21955\,
            I => \N__21952\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__21952\,
            I => \N__21949\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__21949\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1891\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21943\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__21943\,
            I => \pwm_generator_inst.un18_threshold_1_axb_9\
        );

    \I__1889\ : InMux
    port map (
            O => \N__21940\,
            I => \N__21937\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__21937\,
            I => \N__21934\
        );

    \I__1887\ : Span4Mux_v
    port map (
            O => \N__21934\,
            I => \N__21931\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__21931\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1885\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21925\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__21925\,
            I => \pwm_generator_inst.un18_threshold_1_axb_10\
        );

    \I__1883\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21916\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__21916\,
            I => \N__21913\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__21913\,
            I => \pwm_generator_inst.O_11\
        );

    \I__1879\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21907\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__21907\,
            I => \pwm_generator_inst.un18_threshold_1_axb_11\
        );

    \I__1877\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21901\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__21901\,
            I => \N__21898\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__21895\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1873\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__21889\,
            I => \pwm_generator_inst.un18_threshold_1_axb_12\
        );

    \I__1871\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__21880\,
            I => \N__21877\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__21877\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1867\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__21871\,
            I => \pwm_generator_inst.un18_threshold_1_axb_13\
        );

    \I__1865\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21865\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21862\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__21862\,
            I => \N__21859\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__21859\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1861\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21853\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__21853\,
            I => \pwm_generator_inst.un18_threshold_1_axb_0\
        );

    \I__1859\ : InMux
    port map (
            O => \N__21850\,
            I => \N__21847\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21844\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__21844\,
            I => \N__21841\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__21841\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1855\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21835\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__21835\,
            I => \pwm_generator_inst.un18_threshold_1_axb_1\
        );

    \I__1853\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__21829\,
            I => \N__21826\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__21826\,
            I => \N__21823\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__21823\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1849\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__21817\,
            I => \pwm_generator_inst.un18_threshold_1_axb_2\
        );

    \I__1847\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21808\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__21808\,
            I => \N__21805\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__21805\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1843\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__21799\,
            I => \pwm_generator_inst.un18_threshold_1_axb_3\
        );

    \I__1841\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__21787\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1837\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__21781\,
            I => \pwm_generator_inst.un18_threshold_1_axb_4\
        );

    \I__1835\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21772\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__21769\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1831\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21763\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__21763\,
            I => \pwm_generator_inst.un18_threshold_1_axb_5\
        );

    \I__1829\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21757\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__21757\,
            I => \N__21754\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__21754\,
            I => \N__21751\
        );

    \I__1826\ : Sp12to4
    port map (
            O => \N__21751\,
            I => \N__21748\
        );

    \I__1825\ : Span12Mux_s8_h
    port map (
            O => \N__21748\,
            I => \N__21745\
        );

    \I__1824\ : Span12Mux_h
    port map (
            O => \N__21745\,
            I => \N__21742\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__21742\,
            I => \pwm_generator_inst.O_0_1\
        );

    \I__1822\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21736\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__21736\,
            I => \N__21733\
        );

    \I__1820\ : Span4Mux_v
    port map (
            O => \N__21733\,
            I => \N__21730\
        );

    \I__1819\ : Sp12to4
    port map (
            O => \N__21730\,
            I => \N__21727\
        );

    \I__1818\ : Span12Mux_s9_h
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__21721\,
            I => \pwm_generator_inst.O_0_0\
        );

    \I__1815\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__1812\ : Sp12to4
    port map (
            O => \N__21709\,
            I => \N__21706\
        );

    \I__1811\ : Span12Mux_v
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__1810\ : Span12Mux_h
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__1809\ : Span12Mux_v
    port map (
            O => \N__21700\,
            I => \N__21697\
        );

    \I__1808\ : Odrv12
    port map (
            O => \N__21697\,
            I => \pwm_generator_inst.O_0_5\
        );

    \I__1807\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21691\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__21691\,
            I => \N__21688\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__21688\,
            I => \N__21685\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__1803\ : Span12Mux_s6_h
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__1802\ : Span12Mux_h
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__1801\ : Odrv12
    port map (
            O => \N__21676\,
            I => \pwm_generator_inst.O_0_3\
        );

    \I__1800\ : InMux
    port map (
            O => \N__21673\,
            I => \N__21670\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21667\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__21667\,
            I => \N__21664\
        );

    \I__1797\ : Span4Mux_h
    port map (
            O => \N__21664\,
            I => \N__21661\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__21658\,
            I => \N__21655\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__21649\,
            I => \pwm_generator_inst.O_0_4\
        );

    \I__1791\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__1788\ : Sp12to4
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__1787\ : Span12Mux_s7_h
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__1786\ : Span12Mux_h
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__1785\ : Odrv12
    port map (
            O => \N__21628\,
            I => \pwm_generator_inst.O_0_2\
        );

    \I__1784\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__21622\,
            I => \N__21619\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__1780\ : Span12Mux_h
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__1779\ : Span12Mux_h
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__1778\ : Odrv12
    port map (
            O => \N__21607\,
            I => \pwm_generator_inst.O_0_6\
        );

    \I__1777\ : IoInMux
    port map (
            O => \N__21604\,
            I => \N__21601\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__21601\,
            I => \N__21598\
        );

    \I__1775\ : Span4Mux_s3_v
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__1773\ : Sp12to4
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__1772\ : Span12Mux_v
    port map (
            O => \N__21589\,
            I => \N__21586\
        );

    \I__1771\ : Span12Mux_v
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__21583\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1769\ : IoInMux
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21574\
        );

    \I__1767\ : IoSpan4Mux
    port map (
            O => \N__21574\,
            I => \N__21571\
        );

    \I__1766\ : IoSpan4Mux
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__21568\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un22_threshold_1_cry_7\,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_12_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_12_23_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un5_threshold_add_1_cry_7\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un5_threshold_add_1_cry_15\,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un18_threshold_1_cry_7\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un18_threshold_1_cry_15\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un18_threshold_1_cry_23\,
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_4_19_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            carryinitout => \bfn_7_18_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un6_running_cry_30\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_7\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_15\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.counter_cry_23\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un6_running_cry_30\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_7\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_15\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.counter_cry_23\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un6_running_cry_30\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_7\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_15\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.counter_cry_23\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un6_running_cry_30\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\,
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_7\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_15\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.counter_cry_23\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_18_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_7_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_13_20_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21604\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21580\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__30499\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst1.stoper_tr.un2_start_0_g\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29281\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un2_start_0_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__47017\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_163_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__51292\,
            CLKHFEN => \N__51293\,
            CLKHF => clk_12mhz
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21868\,
            in1 => \N__21856\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21838\,
            in2 => \_gnd_net_\,
            in3 => \N__21850\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21832\,
            in1 => \N__21820\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21814\,
            in1 => \N__21802\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21784\,
            in2 => \_gnd_net_\,
            in3 => \N__21796\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21766\,
            in2 => \_gnd_net_\,
            in3 => \N__21778\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22000\,
            in2 => \_gnd_net_\,
            in3 => \N__22012\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21982\,
            in2 => \_gnd_net_\,
            in3 => \N__21994\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21964\,
            in2 => \_gnd_net_\,
            in3 => \N__21976\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21946\,
            in2 => \_gnd_net_\,
            in3 => \N__21958\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21928\,
            in2 => \_gnd_net_\,
            in3 => \N__21940\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21910\,
            in2 => \_gnd_net_\,
            in3 => \N__21922\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21892\,
            in2 => \_gnd_net_\,
            in3 => \N__21904\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21874\,
            in2 => \_gnd_net_\,
            in3 => \N__21886\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22036\,
            in2 => \_gnd_net_\,
            in3 => \N__22048\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22198\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22159\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22264\,
            in2 => \_gnd_net_\,
            in3 => \N__22030\,
            lcout => \pwm_generator_inst.un22_threshold_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22234\,
            in2 => \_gnd_net_\,
            in3 => \N__22027\,
            lcout => \pwm_generator_inst.un18_threshold1_18\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22072\,
            in2 => \_gnd_net_\,
            in3 => \N__22024\,
            lcout => \pwm_generator_inst.un18_threshold1_19\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_18\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22249\,
            in2 => \_gnd_net_\,
            in3 => \N__22021\,
            lcout => \pwm_generator_inst.un18_threshold1_20\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_19\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22066\,
            in2 => \_gnd_net_\,
            in3 => \N__22018\,
            lcout => \pwm_generator_inst.un18_threshold1_21\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_20\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22060\,
            in2 => \_gnd_net_\,
            in3 => \N__22015\,
            lcout => \pwm_generator_inst.un18_threshold1_22\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_21\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22054\,
            in2 => \_gnd_net_\,
            in3 => \N__22084\,
            lcout => \pwm_generator_inst.un18_threshold1_23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_22\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22240\,
            in2 => \_gnd_net_\,
            in3 => \N__22081\,
            lcout => \pwm_generator_inst.un18_threshold1_24\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22255\,
            in2 => \_gnd_net_\,
            in3 => \N__22078\,
            lcout => \pwm_generator_inst.un18_threshold1_25\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un18_threshold_1_cry_24\,
            carryout => \pwm_generator_inst.un18_threshold_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010100110"
        )
    port map (
            in0 => \N__22657\,
            in1 => \N__23393\,
            in2 => \N__23494\,
            in3 => \N__22075\,
            lcout => \pwm_generator_inst.N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23070\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__23509\,
            in1 => \N__23392\,
            in2 => \N__22321\,
            in3 => \N__23523\,
            lcout => \pwm_generator_inst.N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23028\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23295\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23007\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23469\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23457\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23046\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22317\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23343\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22225\,
            in2 => \N__22213\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22189\,
            in2 => \N__22177\,
            in3 => \N__22150\,
            lcout => \pwm_generator_inst.un18_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22147\,
            in2 => \N__22135\,
            in3 => \N__22117\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22114\,
            in2 => \N__22102\,
            in3 => \N__22087\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22504\,
            in2 => \N__22492\,
            in3 => \N__22477\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22474\,
            in2 => \N__22462\,
            in3 => \N__22447\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22444\,
            in2 => \N__22432\,
            in3 => \N__22417\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22414\,
            in2 => \N__22402\,
            in3 => \N__22387\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22384\,
            in2 => \N__22369\,
            in3 => \N__22354\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0\,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22351\,
            in2 => \N__22336\,
            in3 => \N__22300\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22297\,
            in2 => \N__22282\,
            in3 => \N__22267\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22579\,
            in2 => \N__22672\,
            in3 => \N__22648\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22645\,
            in2 => \N__22590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22583\,
            in2 => \N__22633\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22618\,
            in2 => \N__22591\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22587\,
            in2 => \N__22603\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un5_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un5_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22510\,
            in2 => \_gnd_net_\,
            in3 => \N__22606\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__22589\,
            in1 => \N__23121\,
            in2 => \_gnd_net_\,
            in3 => \N__22533\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22588\,
            in2 => \_gnd_net_\,
            in3 => \N__22546\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010010110"
        )
    port map (
            in0 => \N__23086\,
            in1 => \N__23122\,
            in2 => \N__22537\,
            in3 => \N__22534\,
            lcout => \pwm_generator_inst.un5_threshold_add_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51949\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22918\,
            in3 => \N__22885\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50900\,
            in2 => \N__22882\,
            in3 => \N__22849\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22846\,
            in2 => \N__51060\,
            in3 => \N__22807\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22804\,
            in2 => \_gnd_net_\,
            in3 => \N__22777\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22774\,
            in2 => \N__51061\,
            in3 => \N__22738\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22735\,
            in2 => \_gnd_net_\,
            in3 => \N__22708\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22705\,
            in2 => \_gnd_net_\,
            in3 => \N__22675\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28216\,
            in2 => \_gnd_net_\,
            in3 => \N__22984\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0\,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28156\,
            in2 => \_gnd_net_\,
            in3 => \N__22975\,
            lcout => \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28108\,
            in2 => \_gnd_net_\,
            in3 => \N__22966\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28051\,
            in2 => \_gnd_net_\,
            in3 => \N__22957\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28015\,
            in2 => \_gnd_net_\,
            in3 => \N__22948\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27991\,
            in2 => \_gnd_net_\,
            in3 => \N__22939\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27961\,
            in2 => \_gnd_net_\,
            in3 => \N__22930\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27928\,
            in2 => \_gnd_net_\,
            in3 => \N__22921\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28501\,
            in2 => \_gnd_net_\,
            in3 => \N__23143\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28462\,
            in2 => \_gnd_net_\,
            in3 => \N__23134\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28435\,
            in2 => \_gnd_net_\,
            in3 => \N__23125\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28312\,
            in2 => \_gnd_net_\,
            in3 => \N__23107\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__28291\,
            in2 => \N__28414\,
            in3 => \N__23089\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__23266\,
            in1 => \N__23278\,
            in2 => \N__23077\,
            in3 => \N__23383\,
            lcout => \pwm_generator_inst.N_181_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__23253\,
            in1 => \N__23239\,
            in2 => \N__23056\,
            in3 => \N__23384\,
            lcout => \pwm_generator_inst.N_182_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__23215\,
            in1 => \N__23227\,
            in2 => \N__23035\,
            in3 => \N__23385\,
            lcout => \pwm_generator_inst.N_183_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__23179\,
            in2 => \N__23167\,
            in3 => \N__23011\,
            lcout => \pwm_generator_inst.N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__23188\,
            in1 => \N__23202\,
            in2 => \N__23302\,
            in3 => \N__23394\,
            lcout => \pwm_generator_inst.N_184_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23481\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51062\,
            in2 => \N__23412\,
            in3 => \N__23281\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23277\,
            in2 => \N__51289\,
            in3 => \N__23257\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51066\,
            in2 => \N__23254\,
            in3 => \N__23230\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23226\,
            in2 => \N__51290\,
            in3 => \N__23206\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51070\,
            in2 => \N__23203\,
            in3 => \N__23182\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23178\,
            in2 => \N__51291\,
            in3 => \N__23155\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51074\,
            in2 => \N__23524\,
            in3 => \N__23503\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un22_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50989\,
            in2 => \N__23439\,
            in3 => \N__23500\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \pwm_generator_inst.un22_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23497\,
            lcout => \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23387\,
            in1 => \N__23485\,
            in2 => \_gnd_net_\,
            in3 => \N__23470\,
            lcout => \pwm_generator_inst.N_179_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__23458\,
            in1 => \N__23391\,
            in2 => \N__23440\,
            in3 => \N__23425\,
            lcout => \pwm_generator_inst.N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__23419\,
            in1 => \N__23413\,
            in2 => \N__23395\,
            in3 => \N__23344\,
            lcout => \pwm_generator_inst.N_180_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23759\,
            in1 => \N__23323\,
            in2 => \N__23332\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23739\,
            in1 => \N__23308\,
            in2 => \N__23317\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23662\,
            in2 => \N__23677\,
            in3 => \N__23717\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23696\,
            in1 => \N__23641\,
            in2 => \N__23656\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23620\,
            in2 => \N__23635\,
            in3 => \N__23972\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23614\,
            in2 => \N__23608\,
            in3 => \N__23952\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23584\,
            in2 => \N__23599\,
            in3 => \N__23930\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23566\,
            in2 => \N__23578\,
            in3 => \N__23909\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23551\,
            in2 => \N__23560\,
            in3 => \N__23888\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23530\,
            in2 => \N__23545\,
            in3 => \N__23819\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23800\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52609\,
            ce => 'H',
            sr => \N__52268\
        );

    \pwm_generator_inst.counter_RNITBL3_9_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23890\,
            in1 => \N__23821\,
            in2 => \_gnd_net_\,
            in3 => \N__23951\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIRPD2_0_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23760\,
            in2 => \_gnd_net_\,
            in3 => \N__23738\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_2_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__23973\,
            in1 => \N__23697\,
            in2 => \N__23773\,
            in3 => \N__23718\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_6_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23770\,
            in1 => \N__23910\,
            in2 => \N__23764\,
            in3 => \N__23932\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23861\,
            in1 => \N__23761\,
            in2 => \_gnd_net_\,
            in3 => \N__23743\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_1_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23857\,
            in1 => \N__23740\,
            in2 => \_gnd_net_\,
            in3 => \N__23722\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_2_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23862\,
            in1 => \N__23719\,
            in2 => \_gnd_net_\,
            in3 => \N__23701\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_3_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23858\,
            in1 => \N__23698\,
            in2 => \_gnd_net_\,
            in3 => \N__23680\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_4_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23863\,
            in1 => \N__23974\,
            in2 => \_gnd_net_\,
            in3 => \N__23956\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_5_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23859\,
            in1 => \N__23953\,
            in2 => \_gnd_net_\,
            in3 => \N__23935\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_6_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23864\,
            in1 => \N__23931\,
            in2 => \_gnd_net_\,
            in3 => \N__23914\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_7_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23860\,
            in1 => \N__23911\,
            in2 => \_gnd_net_\,
            in3 => \N__23893\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__52601\,
            ce => 'H',
            sr => \N__52266\
        );

    \pwm_generator_inst.counter_8_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23866\,
            in1 => \N__23889\,
            in2 => \_gnd_net_\,
            in3 => \N__23869\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__52594\,
            ce => 'H',
            sr => \N__52269\
        );

    \pwm_generator_inst.counter_9_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__23820\,
            in1 => \N__23865\,
            in2 => \_gnd_net_\,
            in3 => \N__23824\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52594\,
            ce => 'H',
            sr => \N__52269\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__24016\,
            in1 => \N__31810\,
            in2 => \N__31840\,
            in3 => \N__24007\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_16_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52621\,
            ce => \N__36636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__24015\,
            in1 => \N__31809\,
            in2 => \N__31839\,
            in3 => \N__24006\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_17_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25680\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52621\,
            ce => \N__36636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__32047\,
            in1 => \N__32067\,
            in2 => \N__23997\,
            in3 => \N__23983\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_18_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25656\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52621\,
            ce => \N__36636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__32046\,
            in1 => \N__32068\,
            in2 => \N__23998\,
            in3 => \N__23982\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_19_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25788\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52621\,
            ce => \N__36636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28684\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52610\,
            ce => \N__32635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_27_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28636\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52610\,
            ce => \N__32635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_26_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28660\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52610\,
            ce => \N__32635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_24_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52610\,
            ce => \N__32635\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_21_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25768\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52602\,
            ce => \N__36637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__26239\,
            in1 => \N__24049\,
            in2 => \N__26215\,
            in3 => \N__24058\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_16_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25711\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52595\,
            ce => \N__32636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101001101"
        )
    port map (
            in0 => \N__26238\,
            in1 => \N__24048\,
            in2 => \N__26214\,
            in3 => \N__24057\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_17_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25684\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52595\,
            ce => \N__32636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__26161\,
            in1 => \N__26184\,
            in2 => \N__24039\,
            in3 => \N__24025\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_18_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25660\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52595\,
            ce => \N__32636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__26160\,
            in1 => \N__26185\,
            in2 => \N__24040\,
            in3 => \N__24024\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_19_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25792\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52595\,
            ce => \N__32636\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__26458\,
            in1 => \N__24121\,
            in2 => \N__26434\,
            in3 => \N__24109\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101001101"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__24120\,
            in2 => \N__26433\,
            in3 => \N__24108\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__24097\,
            in1 => \N__26374\,
            in2 => \N__26403\,
            in3 => \N__24085\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__24096\,
            in1 => \N__26373\,
            in2 => \N__26404\,
            in3 => \N__24084\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24335\,
            in1 => \N__29828\,
            in2 => \_gnd_net_\,
            in3 => \N__24073\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24370\,
            in1 => \N__29783\,
            in2 => \_gnd_net_\,
            in3 => \N__24070\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24336\,
            in1 => \N__24904\,
            in2 => \_gnd_net_\,
            in3 => \N__24067\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24371\,
            in1 => \N__24882\,
            in2 => \_gnd_net_\,
            in3 => \N__24064\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24337\,
            in1 => \N__25139\,
            in2 => \_gnd_net_\,
            in3 => \N__24061\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24372\,
            in1 => \N__25113\,
            in2 => \_gnd_net_\,
            in3 => \N__24148\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24338\,
            in1 => \N__25089\,
            in2 => \_gnd_net_\,
            in3 => \N__24145\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24373\,
            in1 => \N__25065\,
            in2 => \_gnd_net_\,
            in3 => \N__24142\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__52656\,
            ce => \N__36565\,
            sr => \N__52211\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24342\,
            in1 => \N__25041\,
            in2 => \_gnd_net_\,
            in3 => \N__24139\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24355\,
            in1 => \N__25020\,
            in2 => \_gnd_net_\,
            in3 => \N__24136\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24339\,
            in1 => \N__24996\,
            in2 => \_gnd_net_\,
            in3 => \N__24133\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24352\,
            in1 => \N__24974\,
            in2 => \_gnd_net_\,
            in3 => \N__24130\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24340\,
            in1 => \N__25329\,
            in2 => \_gnd_net_\,
            in3 => \N__24127\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24353\,
            in1 => \N__25305\,
            in2 => \_gnd_net_\,
            in3 => \N__24124\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24341\,
            in1 => \N__25281\,
            in2 => \_gnd_net_\,
            in3 => \N__24175\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24354\,
            in1 => \N__25257\,
            in2 => \_gnd_net_\,
            in3 => \N__24172\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__52651\,
            ce => \N__36564\,
            sr => \N__52218\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24364\,
            in1 => \N__25233\,
            in2 => \_gnd_net_\,
            in3 => \N__24169\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24360\,
            in1 => \N__25212\,
            in2 => \_gnd_net_\,
            in3 => \N__24166\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24365\,
            in1 => \N__25188\,
            in2 => \_gnd_net_\,
            in3 => \N__24163\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24361\,
            in1 => \N__25166\,
            in2 => \_gnd_net_\,
            in3 => \N__24160\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24366\,
            in1 => \N__25548\,
            in2 => \_gnd_net_\,
            in3 => \N__24157\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24362\,
            in1 => \N__25524\,
            in2 => \_gnd_net_\,
            in3 => \N__24154\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24367\,
            in1 => \N__25500\,
            in2 => \_gnd_net_\,
            in3 => \N__24151\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24363\,
            in1 => \N__25476\,
            in2 => \_gnd_net_\,
            in3 => \N__24205\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__52644\,
            ce => \N__36557\,
            sr => \N__52224\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24356\,
            in1 => \N__25452\,
            in2 => \_gnd_net_\,
            in3 => \N__24202\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__52639\,
            ce => \N__36556\,
            sr => \N__52233\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24368\,
            in1 => \N__25428\,
            in2 => \_gnd_net_\,
            in3 => \N__24199\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__52639\,
            ce => \N__36556\,
            sr => \N__52233\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24357\,
            in1 => \N__25392\,
            in2 => \_gnd_net_\,
            in3 => \N__24196\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__52639\,
            ce => \N__36556\,
            sr => \N__52233\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24369\,
            in1 => \N__25356\,
            in2 => \_gnd_net_\,
            in3 => \N__24193\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__52639\,
            ce => \N__36556\,
            sr => \N__52233\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24358\,
            in1 => \N__25408\,
            in2 => \_gnd_net_\,
            in3 => \N__24190\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__52639\,
            ce => \N__36556\,
            sr => \N__52233\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__25372\,
            in1 => \N__24359\,
            in2 => \_gnd_net_\,
            in3 => \N__24187\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52639\,
            ce => \N__36556\,
            sr => \N__52233\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33752\,
            in1 => \N__24184\,
            in2 => \_gnd_net_\,
            in3 => \N__27106\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24178\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33753\,
            in1 => \N__24235\,
            in2 => \_gnd_net_\,
            in3 => \N__27031\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => \elapsed_time_ns_1_RNI7IPBB_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24229\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33750\,
            in1 => \N__25612\,
            in2 => \_gnd_net_\,
            in3 => \N__26956\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33749\,
            in1 => \N__24226\,
            in2 => \_gnd_net_\,
            in3 => \N__29628\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => \elapsed_time_ns_1_RNIJI91B_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24220\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24217\,
            in1 => \N__27018\,
            in2 => \_gnd_net_\,
            in3 => \N__33751\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36699\,
            in2 => \_gnd_net_\,
            in3 => \N__36740\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52626\,
            ce => \N__32596\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26914\,
            in1 => \N__25570\,
            in2 => \_gnd_net_\,
            in3 => \N__33776\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24216\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26998\,
            in1 => \N__25591\,
            in2 => \_gnd_net_\,
            in3 => \N__33777\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36502\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24244\,
            in1 => \N__27310\,
            in2 => \_gnd_net_\,
            in3 => \N__33778\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => \elapsed_time_ns_1_RNI6GOBB_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24238\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30090\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30120\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30264\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30105\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30057\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_15_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34227\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_14_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34281\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30042\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52611\,
            ce => \N__32615\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_2_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30028\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34107\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_13_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30069\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34167\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34194\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34137\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_12_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34254\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32754\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52603\,
            ce => \N__32637\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__26109\,
            in1 => \N__24436\,
            in2 => \N__26136\,
            in3 => \N__24445\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32154\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52596\,
            ce => \N__32619\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101001101"
        )
    port map (
            in0 => \N__26110\,
            in1 => \N__24435\,
            in2 => \N__26137\,
            in3 => \N__24444\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25761\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52596\,
            ce => \N__32619\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__26059\,
            in1 => \N__24427\,
            in2 => \N__26089\,
            in3 => \N__24418\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__26058\,
            in1 => \N__24426\,
            in2 => \N__26088\,
            in3 => \N__24417\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32679\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52596\,
            ce => \N__32619\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24409\,
            in2 => \N__24400\,
            in3 => \N__25893\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24379\,
            in2 => \N__24391\,
            in3 => \N__25881\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24583\,
            in2 => \N__24595\,
            in3 => \N__25866\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24565\,
            in2 => \N__24577\,
            in3 => \N__25851\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24559\,
            in2 => \N__24544\,
            in3 => \N__25836\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24523\,
            in2 => \N__24535\,
            in3 => \N__25821\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24517\,
            in2 => \N__24508\,
            in3 => \N__25806\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26034\,
            in1 => \N__24487\,
            in2 => \N__24499\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26019\,
            in1 => \N__24481\,
            in2 => \N__24472\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_7_18_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26004\,
            in1 => \N__24451\,
            in2 => \N__24463\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24760\,
            in2 => \N__24751\,
            in3 => \N__25989\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24730\,
            in2 => \N__24742\,
            in3 => \N__25974\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24724\,
            in2 => \N__24715\,
            in3 => \N__25959\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24706\,
            in2 => \N__24697\,
            in3 => \N__25944\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24673\,
            in2 => \N__24685\,
            in3 => \N__25929\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24667\,
            in2 => \N__24658\,
            in3 => \N__26253\,
            lcout => \phase_controller_inst2.stoper_tr.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24649\,
            in2 => \N__24637\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24622\,
            in2 => \N__24610\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24865\,
            in2 => \N__24856\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24844\,
            in2 => \N__24832\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24820\,
            in2 => \N__24811\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24799\,
            in2 => \N__24790\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24937\,
            in2 => \N__24946\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24952\,
            in2 => \N__24772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un6_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24775\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__32658\,
            in1 => \N__26289\,
            in2 => \_gnd_net_\,
            in3 => \N__26309\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__26310\,
            in1 => \N__26288\,
            in2 => \_gnd_net_\,
            in3 => \N__32659\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__32656\,
            in1 => \N__26327\,
            in2 => \_gnd_net_\,
            in3 => \N__26348\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__26328\,
            in1 => \N__26349\,
            in2 => \_gnd_net_\,
            in3 => \N__32657\,
            lcout => \phase_controller_inst2.stoper_tr.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32556\,
            in2 => \_gnd_net_\,
            in3 => \N__29220\,
            lcout => \phase_controller_inst2.stoper_tr.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24931\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29269\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52652\,
            ce => 'H',
            sr => \N__52199\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24902\,
            in2 => \N__29835\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24881\,
            in2 => \N__29790\,
            in3 => \N__24907\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24903\,
            in2 => \N__25140\,
            in3 => \N__24889\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25112\,
            in2 => \N__24886\,
            in3 => \N__25144\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25088\,
            in2 => \N__25141\,
            in3 => \N__25120\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25064\,
            in2 => \N__25117\,
            in3 => \N__25096\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25040\,
            in2 => \N__25093\,
            in3 => \N__25072\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25019\,
            in2 => \N__25069\,
            in3 => \N__25048\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__52645\,
            ce => \N__36478\,
            sr => \N__52212\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24995\,
            in2 => \N__25045\,
            in3 => \N__25024\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25021\,
            in2 => \N__24975\,
            in3 => \N__25003\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25328\,
            in2 => \N__25000\,
            in3 => \N__24979\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25304\,
            in2 => \N__24976\,
            in3 => \N__24955\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25280\,
            in2 => \N__25333\,
            in3 => \N__25312\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25256\,
            in2 => \N__25309\,
            in3 => \N__25288\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25232\,
            in2 => \N__25285\,
            in3 => \N__25264\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25211\,
            in2 => \N__25261\,
            in3 => \N__25240\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__52640\,
            ce => \N__36477\,
            sr => \N__52219\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25187\,
            in2 => \N__25237\,
            in3 => \N__25216\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25213\,
            in2 => \N__25167\,
            in3 => \N__25195\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25547\,
            in2 => \N__25192\,
            in3 => \N__25171\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25523\,
            in2 => \N__25168\,
            in3 => \N__25147\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25499\,
            in2 => \N__25552\,
            in3 => \N__25531\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25475\,
            in2 => \N__25528\,
            in3 => \N__25507\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25451\,
            in2 => \N__25504\,
            in3 => \N__25483\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25427\,
            in2 => \N__25480\,
            in3 => \N__25459\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__52633\,
            ce => \N__36476\,
            sr => \N__52225\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25391\,
            in2 => \N__25456\,
            in3 => \N__25435\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__52627\,
            ce => \N__36475\,
            sr => \N__52234\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25355\,
            in2 => \N__25432\,
            in3 => \N__25411\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__52627\,
            ce => \N__36475\,
            sr => \N__52234\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25407\,
            in2 => \N__25396\,
            in3 => \N__25375\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__52627\,
            ce => \N__36475\,
            sr => \N__52234\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25371\,
            in2 => \N__25360\,
            in3 => \N__25339\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__52627\,
            ce => \N__36475\,
            sr => \N__52234\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25336\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52627\,
            ce => \N__36475\,
            sr => \N__52234\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25611\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33772\,
            in1 => \N__25600\,
            in2 => \_gnd_net_\,
            in3 => \N__27094\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25594\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25579\,
            in1 => \N__26941\,
            in2 => \_gnd_net_\,
            in3 => \N__33771\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => \elapsed_time_ns_1_RNILK91B_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25573\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25569\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33796\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36691\,
            in1 => \N__25558\,
            in2 => \N__36742\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27268\,
            in1 => \N__27264\,
            in2 => \N__51471\,
            in3 => \N__25639\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_1,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27238\,
            in1 => \N__27231\,
            in2 => \N__51495\,
            in3 => \N__25636\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_2,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27213\,
            in1 => \N__27214\,
            in2 => \N__51472\,
            in3 => \N__25633\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_3,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27181\,
            in1 => \N__27177\,
            in2 => \N__51496\,
            in3 => \N__25630\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_4,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27157\,
            in1 => \N__27156\,
            in2 => \N__51473\,
            in3 => \N__25627\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_5,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27513\,
            in1 => \N__27517\,
            in2 => \N__51497\,
            in3 => \N__25624\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_6,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27490\,
            in1 => \N__27489\,
            in2 => \N__51474\,
            in3 => \N__25621\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_7,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27475\,
            in1 => \N__27474\,
            in2 => \N__51469\,
            in3 => \N__25618\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_8,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27445\,
            in1 => \N__27441\,
            in2 => \N__51466\,
            in3 => \N__25615\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_9,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27421\,
            in1 => \N__27417\,
            in2 => \N__51470\,
            in3 => \N__25729\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_10,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27390\,
            in1 => \N__27391\,
            in2 => \N__51463\,
            in3 => \N__25726\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_11,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27364\,
            in1 => \N__27360\,
            in2 => \N__51467\,
            in3 => \N__25723\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_12,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27330\,
            in1 => \N__27331\,
            in2 => \N__51464\,
            in3 => \N__25720\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_13,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27724\,
            in1 => \N__27723\,
            in2 => \N__51468\,
            in3 => \N__25717\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_14,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27700\,
            in1 => \N__27699\,
            in2 => \N__51465\,
            in3 => \N__25714\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_15,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27676\,
            in1 => \N__27675\,
            in2 => \N__51298\,
            in3 => \N__25687\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_16,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27655\,
            in1 => \N__27651\,
            in2 => \N__51373\,
            in3 => \N__25663\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_17,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27625\,
            in1 => \N__27621\,
            in2 => \N__51299\,
            in3 => \N__25642\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_18,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27600\,
            in1 => \N__27601\,
            in2 => \N__51374\,
            in3 => \N__25774\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_19,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27565\,
            in1 => \N__27561\,
            in2 => \N__51300\,
            in3 => \N__25771\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_20,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27543\,
            in1 => \N__27544\,
            in2 => \N__51375\,
            in3 => \N__25750\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_21,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27910\,
            in1 => \N__27909\,
            in2 => \N__51301\,
            in3 => \N__25747\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_22,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27886\,
            in1 => \N__27885\,
            in2 => \N__51376\,
            in3 => \N__25744\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_23,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27859\,
            in1 => \N__27858\,
            in2 => \N__51294\,
            in3 => \N__25741\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_24,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27838\,
            in1 => \N__27834\,
            in2 => \N__51296\,
            in3 => \N__25738\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_25,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27802\,
            in1 => \N__27798\,
            in2 => \N__51295\,
            in3 => \N__25735\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_26,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27777\,
            in1 => \N__27778\,
            in2 => \N__51297\,
            in3 => \N__25732\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_27,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25915\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.counter_0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32503\,
            in1 => \N__25894\,
            in2 => \N__25912\,
            in3 => \N__25911\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_0\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_1_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32490\,
            in1 => \N__25882\,
            in2 => \_gnd_net_\,
            in3 => \N__25870\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_1\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_2_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32504\,
            in1 => \N__25867\,
            in2 => \_gnd_net_\,
            in3 => \N__25855\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_2\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_3_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32491\,
            in1 => \N__25852\,
            in2 => \_gnd_net_\,
            in3 => \N__25840\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_3\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_4_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32505\,
            in1 => \N__25837\,
            in2 => \_gnd_net_\,
            in3 => \N__25825\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_4\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_5_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32492\,
            in1 => \N__25822\,
            in2 => \_gnd_net_\,
            in3 => \N__25810\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_5\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_6_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32506\,
            in1 => \N__25807\,
            in2 => \_gnd_net_\,
            in3 => \N__25795\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_6\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_7_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32493\,
            in1 => \N__26035\,
            in2 => \_gnd_net_\,
            in3 => \N__26023\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_7\,
            clk => \N__52584\,
            ce => \N__26269\,
            sr => \N__52251\
        );

    \phase_controller_inst2.stoper_tr.counter_8_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32489\,
            in1 => \N__26020\,
            in2 => \_gnd_net_\,
            in3 => \N__26008\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_8\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_9_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32499\,
            in1 => \N__26005\,
            in2 => \_gnd_net_\,
            in3 => \N__25993\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_9\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_10_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32486\,
            in1 => \N__25990\,
            in2 => \_gnd_net_\,
            in3 => \N__25978\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_10\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_11_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32500\,
            in1 => \N__25975\,
            in2 => \_gnd_net_\,
            in3 => \N__25963\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_11\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_12_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32487\,
            in1 => \N__25960\,
            in2 => \_gnd_net_\,
            in3 => \N__25948\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_12\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_13_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32501\,
            in1 => \N__25945\,
            in2 => \_gnd_net_\,
            in3 => \N__25933\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_13\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_14_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32488\,
            in1 => \N__25930\,
            in2 => \_gnd_net_\,
            in3 => \N__25918\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_14\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_15_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32502\,
            in1 => \N__26254\,
            in2 => \_gnd_net_\,
            in3 => \N__26242\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_15\,
            clk => \N__52578\,
            ce => \N__26270\,
            sr => \N__52256\
        );

    \phase_controller_inst2.stoper_tr.counter_16_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32478\,
            in1 => \N__26232\,
            in2 => \_gnd_net_\,
            in3 => \N__26218\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_16\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_17_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32482\,
            in1 => \N__26202\,
            in2 => \_gnd_net_\,
            in3 => \N__26188\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_17\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_18_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32479\,
            in1 => \N__26178\,
            in2 => \_gnd_net_\,
            in3 => \N__26164\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_18\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_19_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32483\,
            in1 => \N__26154\,
            in2 => \_gnd_net_\,
            in3 => \N__26140\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_19\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_20_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32480\,
            in1 => \N__26129\,
            in2 => \_gnd_net_\,
            in3 => \N__26113\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_20\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_21_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32484\,
            in1 => \N__26108\,
            in2 => \_gnd_net_\,
            in3 => \N__26092\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_21\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_22_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32481\,
            in1 => \N__26076\,
            in2 => \_gnd_net_\,
            in3 => \N__26062\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_22\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_23_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32485\,
            in1 => \N__26052\,
            in2 => \_gnd_net_\,
            in3 => \N__26038\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_23\,
            clk => \N__52573\,
            ce => \N__26271\,
            sr => \N__52260\
        );

    \phase_controller_inst2.stoper_tr.counter_24_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32494\,
            in1 => \N__26451\,
            in2 => \_gnd_net_\,
            in3 => \N__26437\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_24\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_25_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32507\,
            in1 => \N__26421\,
            in2 => \_gnd_net_\,
            in3 => \N__26407\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_25\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_26_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32495\,
            in1 => \N__26391\,
            in2 => \_gnd_net_\,
            in3 => \N__26377\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_26\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_27_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32508\,
            in1 => \N__26367\,
            in2 => \_gnd_net_\,
            in3 => \N__26353\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_27\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_28_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32496\,
            in1 => \N__26350\,
            in2 => \_gnd_net_\,
            in3 => \N__26332\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_28\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_29_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32509\,
            in1 => \N__26329\,
            in2 => \_gnd_net_\,
            in3 => \N__26314\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_29\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_30_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32497\,
            in1 => \N__26311\,
            in2 => \_gnd_net_\,
            in3 => \N__26296\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.counter_cry_29\,
            carryout => \phase_controller_inst2.stoper_tr.counter_cry_30\,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \phase_controller_inst2.stoper_tr.counter_31_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26290\,
            in1 => \N__32498\,
            in2 => \_gnd_net_\,
            in3 => \N__26293\,
            lcout => \phase_controller_inst2.stoper_tr.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52567\,
            ce => \N__26272\,
            sr => \N__52262\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26701\,
            in2 => \N__26683\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26662\,
            in2 => \N__26647\,
            in3 => \N__26629\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26626\,
            in2 => \N__26611\,
            in3 => \N__26584\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26581\,
            in2 => \N__26563\,
            in3 => \N__26545\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26542\,
            in2 => \N__30764\,
            in3 => \N__26524\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26521\,
            in2 => \N__30766\,
            in3 => \N__26503\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26500\,
            in2 => \N__30765\,
            in3 => \N__26482\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26479\,
            in2 => \N__30767\,
            in3 => \N__26461\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26848\,
            in2 => \N__30768\,
            in3 => \N__26830\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26827\,
            in2 => \N__30772\,
            in3 => \N__26812\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26809\,
            in2 => \N__30769\,
            in3 => \N__26791\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26788\,
            in2 => \N__30773\,
            in3 => \N__26770\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26767\,
            in2 => \N__30770\,
            in3 => \N__26749\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26746\,
            in2 => \N__30774\,
            in3 => \N__26728\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26725\,
            in2 => \N__30771\,
            in3 => \N__26707\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26704\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52290\,
            in1 => \N__34440\,
            in2 => \_gnd_net_\,
            in3 => \N__34395\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52646\,
            ce => 'H',
            sr => \N__52195\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__26870\,
            in1 => \N__34351\,
            in2 => \N__30955\,
            in3 => \N__29467\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52646\,
            ce => 'H',
            sr => \N__52195\
        );

    \phase_controller_inst2.start_timer_tr_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__29441\,
            in1 => \N__26854\,
            in2 => \N__29409\,
            in3 => \N__29268\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52646\,
            ce => 'H',
            sr => \N__52195\
        );

    \phase_controller_inst2.state_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__26895\,
            in1 => \N__29442\,
            in2 => \N__26878\,
            in3 => \N__29404\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52646\,
            ce => 'H',
            sr => \N__52195\
        );

    \phase_controller_inst2.start_timer_hc_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111100000"
        )
    port map (
            in0 => \N__29375\,
            in1 => \N__26894\,
            in2 => \N__29331\,
            in3 => \N__34435\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52646\,
            ce => 'H',
            sr => \N__52195\
        );

    \phase_controller_inst2.state_2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__26896\,
            in1 => \N__29376\,
            in2 => \N__26877\,
            in3 => \N__29327\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52646\,
            ce => 'H',
            sr => \N__52195\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52292\,
            in1 => \N__29267\,
            in2 => \_gnd_net_\,
            in3 => \N__32537\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26893\,
            in2 => \_gnd_net_\,
            in3 => \N__26869\,
            lcout => \phase_controller_inst2.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29697\,
            in2 => \_gnd_net_\,
            in3 => \N__27054\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26967\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__29466\,
            in1 => \_gnd_net_\,
            in2 => \N__34396\,
            in3 => \N__34430\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29850\,
            in1 => \N__29715\,
            in2 => \N__29812\,
            in3 => \N__29767\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33767\,
            in1 => \N__27744\,
            in2 => \_gnd_net_\,
            in3 => \N__27079\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33709\,
            in1 => \N__27136\,
            in2 => \_gnd_net_\,
            in3 => \N__26923\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26976\,
            in1 => \N__27126\,
            in2 => \N__26997\,
            in3 => \N__29535\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27292\,
            in1 => \N__27004\,
            in2 => \N__26980\,
            in3 => \N__27064\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26977\,
            in1 => \N__33710\,
            in2 => \_gnd_net_\,
            in3 => \N__26968\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29511\,
            in1 => \N__26952\,
            in2 => \N__26940\,
            in3 => \N__26922\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26910\,
            in2 => \N__26899\,
            in3 => \N__33843\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27135\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33693\,
            in1 => \N__27115\,
            in2 => \_gnd_net_\,
            in3 => \N__27127\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27109\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27105\,
            in1 => \N__27090\,
            in2 => \N__29988\,
            in3 => \N__27075\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27043\,
            in1 => \N__33691\,
            in2 => \_gnd_net_\,
            in3 => \N__27058\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => \elapsed_time_ns_1_RNIHG91B_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27034\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29598\,
            in1 => \N__36690\,
            in2 => \_gnd_net_\,
            in3 => \N__33692\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27030\,
            in1 => \N__30003\,
            in2 => \N__27019\,
            in3 => \N__33603\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29664\,
            in1 => \N__27303\,
            in2 => \N__29880\,
            in3 => \N__33807\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29566\,
            in1 => \N__36677\,
            in2 => \N__27286\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27277\,
            in2 => \_gnd_net_\,
            in3 => \N__29751\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29728\,
            in2 => \_gnd_net_\,
            in3 => \N__27271\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29959\,
            in2 => \_gnd_net_\,
            in3 => \N__27247\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27244\,
            in2 => \_gnd_net_\,
            in3 => \N__27217\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29677\,
            in2 => \_gnd_net_\,
            in3 => \N__27193\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27190\,
            in2 => \_gnd_net_\,
            in3 => \N__27160\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29908\,
            in2 => \_gnd_net_\,
            in3 => \N__27139\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27523\,
            in2 => \_gnd_net_\,
            in3 => \N__27499\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27496\,
            in2 => \_gnd_net_\,
            in3 => \N__27478\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29491\,
            in2 => \_gnd_net_\,
            in3 => \N__27457\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27454\,
            in2 => \_gnd_net_\,
            in3 => \N__27424\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33823\,
            in2 => \_gnd_net_\,
            in3 => \N__27400\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27397\,
            in2 => \_gnd_net_\,
            in3 => \N__27373\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27370\,
            in2 => \_gnd_net_\,
            in3 => \N__27343\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27340\,
            in2 => \_gnd_net_\,
            in3 => \N__27313\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29551\,
            in2 => \_gnd_net_\,
            in3 => \N__27712\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27709\,
            in2 => \_gnd_net_\,
            in3 => \N__27688\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27685\,
            in2 => \_gnd_net_\,
            in3 => \N__27658\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30148\,
            in2 => \_gnd_net_\,
            in3 => \N__27634\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27631\,
            in2 => \_gnd_net_\,
            in3 => \N__27604\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29890\,
            in2 => \_gnd_net_\,
            in3 => \N__27580\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27577\,
            in2 => \_gnd_net_\,
            in3 => \N__27547\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29941\,
            in2 => \_gnd_net_\,
            in3 => \N__27526\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30130\,
            in2 => \_gnd_net_\,
            in3 => \N__27898\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27895\,
            in2 => \_gnd_net_\,
            in3 => \N__27874\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27871\,
            in2 => \_gnd_net_\,
            in3 => \N__27841\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27730\,
            in2 => \_gnd_net_\,
            in3 => \N__27817\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27814\,
            in2 => \_gnd_net_\,
            in3 => \N__27781\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33583\,
            in2 => \_gnd_net_\,
            in3 => \N__27760\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29\,
            carryout => \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__36692\,
            in1 => \N__27757\,
            in2 => \_gnd_net_\,
            in3 => \N__27748\,
            lcout => phase_controller_inst1_stoper_tr_target_ticks_1_i_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27745\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28249\,
            in2 => \N__28237\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28195\,
            in2 => \N__28180\,
            in3 => \N__28144\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28141\,
            in2 => \N__28123\,
            in3 => \N__28087\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28084\,
            in2 => \N__28066\,
            in3 => \N__28036\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28388\,
            in2 => \N__28033\,
            in3 => \N__28003\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28000\,
            in2 => \N__28409\,
            in3 => \N__27973\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27970\,
            in2 => \N__28411\,
            in3 => \N__27943\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27940\,
            in2 => \N__28410\,
            in3 => \N__28516\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28513\,
            in2 => \N__28412\,
            in3 => \N__28483\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28401\,
            in2 => \N__28480\,
            in3 => \N__28450\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28447\,
            in2 => \N__28413\,
            in3 => \N__28417\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28405\,
            in2 => \N__28330\,
            in3 => \N__28297\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28294\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100010000"
        )
    port map (
            in0 => \N__31990\,
            in1 => \N__32014\,
            in2 => \N__28264\,
            in3 => \N__28669\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28275\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52579\,
            ce => \N__36624\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__31989\,
            in1 => \N__32013\,
            in2 => \N__28263\,
            in3 => \N__28668\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28680\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52579\,
            ce => \N__36624\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__28645\,
            in1 => \N__32368\,
            in2 => \N__31965\,
            in3 => \N__28621\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28656\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52579\,
            ce => \N__36624\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28644\,
            in1 => \N__32367\,
            in2 => \N__31966\,
            in3 => \N__28620\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_27_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28632\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52579\,
            ce => \N__36624\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34693\,
            in2 => \N__28612\,
            in3 => \N__32878\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \N__52574\,
            ce => 'H',
            sr => \N__52252\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__32877\,
            in1 => \N__34655\,
            in2 => \N__28588\,
            in3 => \N__28567\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \N__52574\,
            ce => 'H',
            sr => \N__52252\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__32880\,
            in1 => \N__34628\,
            in2 => \N__28564\,
            in3 => \N__28543\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \N__52574\,
            ce => 'H',
            sr => \N__52252\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35089\,
            in2 => \N__28540\,
            in3 => \N__28519\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35052\,
            in2 => \N__28876\,
            in3 => \N__28852\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34998\,
            in2 => \N__28849\,
            in3 => \N__28828\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34945\,
            in2 => \N__28825\,
            in3 => \N__28804\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34909\,
            in2 => \N__28801\,
            in3 => \N__28783\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28780\,
            in2 => \N__34860\,
            in3 => \N__28759\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34822\,
            in2 => \N__28756\,
            in3 => \N__28738\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34770\,
            in2 => \N__28735\,
            in3 => \N__28714\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35424\,
            in2 => \N__28711\,
            in3 => \N__28687\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35362\,
            in2 => \N__29014\,
            in3 => \N__28990\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35299\,
            in2 => \N__28987\,
            in3 => \N__28963\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35265\,
            in2 => \N__28960\,
            in3 => \N__28939\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35202\,
            in2 => \N__28936\,
            in3 => \N__28921\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28918\,
            in2 => \N__37619\,
            in3 => \N__28909\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28906\,
            in2 => \N__35157\,
            in3 => \N__28900\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37667\,
            in2 => \N__28897\,
            in3 => \N__28888\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28885\,
            in2 => \N__37704\,
            in3 => \N__28879\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35685\,
            in2 => \N__29131\,
            in3 => \N__29119\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29116\,
            in2 => \N__37580\,
            in3 => \N__29110\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35652\,
            in2 => \N__29107\,
            in3 => \N__29098\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35612\,
            in2 => \N__29095\,
            in3 => \N__29080\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35577\,
            in2 => \N__29077\,
            in3 => \N__29068\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35547\,
            in2 => \N__29065\,
            in3 => \N__29056\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35504\,
            in2 => \N__29053\,
            in3 => \N__29044\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35462\,
            in2 => \N__29041\,
            in3 => \N__29029\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35932\,
            in2 => \N__29026\,
            in3 => \N__29017\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35898\,
            in2 => \N__29209\,
            in3 => \N__29200\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_er_31_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35829\,
            in1 => \N__29197\,
            in2 => \N__30670\,
            in3 => \N__29191\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52557\,
            ce => \N__32924\,
            sr => \N__52263\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35817\,
            in1 => \N__32917\,
            in2 => \_gnd_net_\,
            in3 => \N__29188\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52553\,
            ce => 'H',
            sr => \N__52264\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32916\,
            in1 => \N__35820\,
            in2 => \_gnd_net_\,
            in3 => \N__29182\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52553\,
            ce => 'H',
            sr => \N__52264\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35818\,
            in1 => \N__32918\,
            in2 => \_gnd_net_\,
            in3 => \N__29176\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52553\,
            ce => 'H',
            sr => \N__52264\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32915\,
            in1 => \N__35819\,
            in2 => \_gnd_net_\,
            in3 => \N__29170\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52553\,
            ce => 'H',
            sr => \N__52264\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32925\,
            in1 => \N__35856\,
            in2 => \_gnd_net_\,
            in3 => \N__29161\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52548\,
            ce => 'H',
            sr => \N__52267\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35855\,
            in1 => \N__29152\,
            in2 => \_gnd_net_\,
            in3 => \N__32926\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52548\,
            ce => 'H',
            sr => \N__52267\
        );

    \phase_controller_inst2.S1_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29335\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52545\,
            ce => 'H',
            sr => \N__52270\
        );

    \phase_controller_inst2.S2_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29419\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52540\,
            ce => 'H',
            sr => \N__52271\
        );

    \phase_controller_inst2.stoper_hc.running_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011101110"
        )
    port map (
            in0 => \N__34434\,
            in1 => \N__29465\,
            in2 => \N__30954\,
            in3 => \N__34386\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52641\,
            ce => 'H',
            sr => \N__52178\
        );

    \phase_controller_inst2.state_0_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__29298\,
            in1 => \N__29446\,
            in2 => \N__29353\,
            in3 => \N__29405\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52641\,
            ce => 'H',
            sr => \N__52178\
        );

    \phase_controller_inst2.state_RNO_0_3_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__29380\,
            in1 => \N__29323\,
            in2 => \N__29299\,
            in3 => \N__29349\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.state_ns_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__34008\,
            in1 => \N__34063\,
            in2 => \N__29338\,
            in3 => \N__34084\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52635\,
            ce => 'H',
            sr => \N__52187\
        );

    \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29265\,
            in2 => \_gnd_net_\,
            in3 => \N__32545\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_tr.un4_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__29653\,
            in1 => \N__29297\,
            in2 => \N__29302\,
            in3 => \N__29238\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52635\,
            ce => 'H',
            sr => \N__52187\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__29651\,
            in1 => \N__29264\,
            in2 => \_gnd_net_\,
            in3 => \N__32544\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__29266\,
            in1 => \N__29652\,
            in2 => \N__32555\,
            in3 => \N__29239\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52635\,
            ce => 'H',
            sr => \N__52187\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_25_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41143\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52629\,
            ce => \N__41915\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__29934\,
            in1 => \N__29638\,
            in2 => \N__29632\,
            in3 => \N__29608\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__29602\,
            in1 => \N__29584\,
            in2 => \N__29578\,
            in3 => \N__29575\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29808\,
            in2 => \N__29569\,
            in3 => \N__29565\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29523\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29524\,
            in1 => \_gnd_net_\,
            in2 => \N__33727\,
            in3 => \N__29539\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29500\,
            in1 => \N__29515\,
            in2 => \_gnd_net_\,
            in3 => \N__33682\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => \elapsed_time_ns_1_RNIU7OBB_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29494\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29740\,
            in1 => \N__29857\,
            in2 => \_gnd_net_\,
            in3 => \N__33681\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29839\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52613\,
            ce => \N__36462\,
            sr => \N__52206\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29794\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52613\,
            ce => \N__36462\,
            sr => \N__52206\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29752\,
            in1 => \N__33694\,
            in2 => \_gnd_net_\,
            in3 => \N__29766\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29739\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33695\,
            in1 => \N__29971\,
            in2 => \_gnd_net_\,
            in3 => \N__29722\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29704\,
            in1 => \N__29686\,
            in2 => \_gnd_net_\,
            in3 => \N__33723\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => \elapsed_time_ns_1_RNIIH91B_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29680\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29902\,
            in1 => \N__29671\,
            in2 => \_gnd_net_\,
            in3 => \N__33724\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33725\,
            in1 => \N__29953\,
            in2 => \_gnd_net_\,
            in3 => \N__30010\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30142\,
            in1 => \N__33726\,
            in2 => \_gnd_net_\,
            in3 => \N__29992\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29970\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29952\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29935\,
            in1 => \N__29917\,
            in2 => \_gnd_net_\,
            in3 => \N__33728\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => \elapsed_time_ns_1_RNIKJ91B_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29911\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29901\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29863\,
            in1 => \N__29884\,
            in2 => \_gnd_net_\,
            in3 => \N__33729\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30151\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30141\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_6_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30106\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_5_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30091\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_13_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30076\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_7_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30058\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_4_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30043\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30024\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_3_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30265\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52590\,
            ce => \N__36617\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36649\,
            in2 => \N__30250\,
            in3 => \N__31425\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30241\,
            in2 => \N__30235\,
            in3 => \N__31785\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30217\,
            in2 => \N__30226\,
            in3 => \N__31770\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30211\,
            in2 => \N__30205\,
            in3 => \N__31755\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30196\,
            in2 => \N__30190\,
            in3 => \N__31740\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31726\,
            in1 => \N__30181\,
            in2 => \N__30175\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30166\,
            in2 => \N__30160\,
            in3 => \N__31707\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30358\,
            in2 => \N__30352\,
            in3 => \N__31693\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31674\,
            in1 => \N__30340\,
            in2 => \N__34156\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34123\,
            in2 => \N__30334\,
            in3 => \N__31659\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30325\,
            in2 => \N__34096\,
            in3 => \N__31936\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34183\,
            in2 => \N__30319\,
            in3 => \N__31914\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34243\,
            in2 => \N__30310\,
            in3 => \N__31899\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30301\,
            in2 => \N__30292\,
            in3 => \N__31884\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34270\,
            in2 => \N__30283\,
            in3 => \N__31869\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34213\,
            in2 => \N__30274\,
            in3 => \N__31854\,
            lcout => \phase_controller_inst1.stoper_tr.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30454\,
            in2 => \N__30439\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30421\,
            in2 => \N__30406\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32080\,
            in2 => \N__32173\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32692\,
            in2 => \N__32770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30388\,
            in2 => \N__30382\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30373\,
            in2 => \N__30367\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34591\,
            in2 => \N__34528\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34456\,
            in2 => \N__34516\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un6_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30502\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34315\,
            in1 => \N__36781\,
            in2 => \_gnd_net_\,
            in3 => \N__36816\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36815\,
            in2 => \_gnd_net_\,
            in3 => \N__34326\,
            lcout => \phase_controller_inst1.stoper_tr.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35863\,
            in1 => \N__30478\,
            in2 => \_gnd_net_\,
            in3 => \N__32898\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52563\,
            ce => 'H',
            sr => \N__52245\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__35864\,
            in1 => \N__30472\,
            in2 => \_gnd_net_\,
            in3 => \N__32899\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52563\,
            ce => 'H',
            sr => \N__52245\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__30550\,
            in1 => \N__35094\,
            in2 => \N__34920\,
            in3 => \N__34629\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__33040\,
            in1 => \N__30526\,
            in2 => \N__30466\,
            in3 => \N__32962\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30463\,
            in1 => \_gnd_net_\,
            in2 => \N__30457\,
            in3 => \N__35865\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52563\,
            ce => 'H',
            sr => \N__52245\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34950\,
            in1 => \N__34997\,
            in2 => \N__35051\,
            in3 => \N__34859\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__30544\,
            in1 => \N__35860\,
            in2 => \_gnd_net_\,
            in3 => \N__32881\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52559\,
            ce => 'H',
            sr => \N__52247\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__35859\,
            in1 => \N__32879\,
            in2 => \_gnd_net_\,
            in3 => \N__30538\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52559\,
            ce => 'H',
            sr => \N__52247\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__30532\,
            in1 => \N__35861\,
            in2 => \_gnd_net_\,
            in3 => \N__32882\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52559\,
            ce => 'H',
            sr => \N__52247\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35858\,
            in1 => \N__35150\,
            in2 => \_gnd_net_\,
            in3 => \N__32932\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__34627\,
            in1 => \N__34656\,
            in2 => \N__34701\,
            in3 => \N__35090\,
            lcout => \current_shift_inst.PI_CTRL.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34697\,
            in2 => \_gnd_net_\,
            in3 => \N__34729\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52559\,
            ce => 'H',
            sr => \N__52247\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35822\,
            in1 => \N__30520\,
            in2 => \_gnd_net_\,
            in3 => \N__32905\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32902\,
            in1 => \N__35826\,
            in2 => \_gnd_net_\,
            in3 => \N__30514\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32900\,
            in1 => \N__35825\,
            in2 => \_gnd_net_\,
            in3 => \N__30508\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__35824\,
            in1 => \N__30607\,
            in2 => \_gnd_net_\,
            in3 => \N__32906\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32901\,
            in1 => \N__30598\,
            in2 => \_gnd_net_\,
            in3 => \N__35828\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35823\,
            in1 => \N__32904\,
            in2 => \_gnd_net_\,
            in3 => \N__30592\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32903\,
            in1 => \N__35827\,
            in2 => \_gnd_net_\,
            in3 => \N__30586\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52555\,
            ce => 'H',
            sr => \N__52253\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32907\,
            in1 => \N__35814\,
            in2 => \_gnd_net_\,
            in3 => \N__30580\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52550\,
            ce => 'H',
            sr => \N__52257\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35811\,
            in1 => \N__32910\,
            in2 => \_gnd_net_\,
            in3 => \N__30574\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52550\,
            ce => 'H',
            sr => \N__52257\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32909\,
            in1 => \N__35816\,
            in2 => \_gnd_net_\,
            in3 => \N__30568\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52550\,
            ce => 'H',
            sr => \N__52257\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35813\,
            in1 => \N__32912\,
            in2 => \_gnd_net_\,
            in3 => \N__30562\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52550\,
            ce => 'H',
            sr => \N__52257\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32908\,
            in1 => \N__35815\,
            in2 => \_gnd_net_\,
            in3 => \N__30556\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52550\,
            ce => 'H',
            sr => \N__52257\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35812\,
            in1 => \N__32911\,
            in2 => \_gnd_net_\,
            in3 => \N__30808\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52550\,
            ce => 'H',
            sr => \N__52257\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35821\,
            in1 => \N__30802\,
            in2 => \_gnd_net_\,
            in3 => \N__32914\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52547\,
            ce => 'H',
            sr => \N__52261\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35461\,
            in1 => \N__35503\,
            in2 => \N__35413\,
            in3 => \N__35897\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30793\,
            in2 => \_gnd_net_\,
            in3 => \N__30775\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31102\,
            in1 => \N__41965\,
            in2 => \N__30658\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33298\,
            in2 => \N__30649\,
            in3 => \N__31087\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33004\,
            in2 => \N__30640\,
            in3 => \N__31066\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32998\,
            in2 => \N__30628\,
            in3 => \N__31048\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33088\,
            in2 => \N__30619\,
            in3 => \N__31024\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31006\,
            in1 => \N__32992\,
            in2 => \N__30877\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30988\,
            in1 => \N__33094\,
            in2 => \N__30868\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33100\,
            in2 => \N__30859\,
            in3 => \N__31300\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30850\,
            in2 => \N__32986\,
            in3 => \N__31279\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33010\,
            in2 => \N__30844\,
            in3 => \N__31258\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33292\,
            in2 => \N__30835\,
            in3 => \N__31240\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30826\,
            in2 => \N__33076\,
            in3 => \N__31222\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33055\,
            in2 => \N__30820\,
            in3 => \N__31204\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33082\,
            in2 => \N__30907\,
            in3 => \N__31186\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31165\,
            in1 => \N__33067\,
            in2 => \N__30898\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33061\,
            in2 => \N__30886\,
            in3 => \N__31147\,
            lcout => \phase_controller_inst2.stoper_hc.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33286\,
            in2 => \N__33223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30961\,
            in2 => \N__33130\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30967\,
            in2 => \N__31126\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30913\,
            in2 => \N__30922\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33307\,
            in2 => \N__33505\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33493\,
            in2 => \N__33430\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33406\,
            in2 => \N__33364\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33925\,
            in2 => \N__33865\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un6_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30970\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100001010"
        )
    port map (
            in0 => \N__33349\,
            in1 => \N__31402\,
            in2 => \N__31381\,
            in3 => \N__33109\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__33189\,
            in1 => \N__33205\,
            in2 => \N__33166\,
            in3 => \N__33121\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34397\,
            in2 => \_gnd_net_\,
            in3 => \N__30938\,
            lcout => \phase_controller_inst2.stoper_hc.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001110"
        )
    port map (
            in0 => \N__33331\,
            in1 => \N__33340\,
            in2 => \N__31327\,
            in3 => \N__31353\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__33339\,
            in1 => \N__33330\,
            in2 => \N__31354\,
            in3 => \N__31326\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100101011"
        )
    port map (
            in0 => \N__33348\,
            in1 => \N__31401\,
            in2 => \N__31380\,
            in3 => \N__33108\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.counter_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31575\,
            in1 => \N__31101\,
            in2 => \N__31117\,
            in3 => \N__31116\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_0\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31613\,
            in1 => \N__31083\,
            in2 => \_gnd_net_\,
            in3 => \N__31069\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_1\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31576\,
            in1 => \N__31065\,
            in2 => \_gnd_net_\,
            in3 => \N__31051\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_2\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__31614\,
            in1 => \_gnd_net_\,
            in2 => \N__31047\,
            in3 => \N__31027\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_3\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_4_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31577\,
            in1 => \N__31023\,
            in2 => \_gnd_net_\,
            in3 => \N__31009\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_4\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31615\,
            in1 => \N__31005\,
            in2 => \_gnd_net_\,
            in3 => \N__30991\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_5\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_6_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31578\,
            in1 => \N__30987\,
            in2 => \_gnd_net_\,
            in3 => \N__30973\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_6\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_7_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31616\,
            in1 => \N__31296\,
            in2 => \_gnd_net_\,
            in3 => \N__31282\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_7\,
            clk => \N__52614\,
            ce => \N__31490\,
            sr => \N__52191\
        );

    \phase_controller_inst2.stoper_hc.counter_8_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31600\,
            in1 => \N__31275\,
            in2 => \_gnd_net_\,
            in3 => \N__31261\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_8\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_9_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31612\,
            in1 => \N__31257\,
            in2 => \_gnd_net_\,
            in3 => \N__31243\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_9\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_10_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31597\,
            in1 => \N__31239\,
            in2 => \_gnd_net_\,
            in3 => \N__31225\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_10\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_11_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31609\,
            in1 => \N__31221\,
            in2 => \_gnd_net_\,
            in3 => \N__31207\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_11\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_12_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31598\,
            in1 => \N__31203\,
            in2 => \_gnd_net_\,
            in3 => \N__31189\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_12\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_13_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31610\,
            in1 => \N__31182\,
            in2 => \_gnd_net_\,
            in3 => \N__31168\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_13\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_14_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31599\,
            in1 => \N__31164\,
            in2 => \_gnd_net_\,
            in3 => \N__31150\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_14\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_15_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31611\,
            in1 => \N__31143\,
            in2 => \_gnd_net_\,
            in3 => \N__31129\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_15\,
            clk => \N__52605\,
            ce => \N__31489\,
            sr => \N__52196\
        );

    \phase_controller_inst2.stoper_hc.counter_16_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31601\,
            in1 => \N__33237\,
            in2 => \_gnd_net_\,
            in3 => \N__31414\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_16\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_17_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31605\,
            in1 => \N__33264\,
            in2 => \_gnd_net_\,
            in3 => \N__31411\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_17\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_18_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31602\,
            in1 => \N__33152\,
            in2 => \_gnd_net_\,
            in3 => \N__31408\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_18\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_19_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31606\,
            in1 => \N__33185\,
            in2 => \_gnd_net_\,
            in3 => \N__31405\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_19\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_20_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31603\,
            in1 => \N__31400\,
            in2 => \_gnd_net_\,
            in3 => \N__31384\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_20\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_21_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31607\,
            in1 => \N__31373\,
            in2 => \_gnd_net_\,
            in3 => \N__31357\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_21\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_22_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31604\,
            in1 => \N__31344\,
            in2 => \_gnd_net_\,
            in3 => \N__31330\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_22\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_23_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31608\,
            in1 => \N__31317\,
            in2 => \_gnd_net_\,
            in3 => \N__31303\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_23\,
            clk => \N__52598\,
            ce => \N__31491\,
            sr => \N__52207\
        );

    \phase_controller_inst2.stoper_hc.counter_24_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31617\,
            in1 => \N__33521\,
            in2 => \_gnd_net_\,
            in3 => \N__31645\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_24\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_25_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31622\,
            in1 => \N__33560\,
            in2 => \_gnd_net_\,
            in3 => \N__31642\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_25\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_26_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31618\,
            in1 => \N__33444\,
            in2 => \_gnd_net_\,
            in3 => \N__31639\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_26\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_27_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31623\,
            in1 => \N__33473\,
            in2 => \_gnd_net_\,
            in3 => \N__31636\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_27\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_28_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31619\,
            in1 => \N__33379\,
            in2 => \_gnd_net_\,
            in3 => \N__31633\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_28\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_29_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31624\,
            in1 => \N__33394\,
            in2 => \_gnd_net_\,
            in3 => \N__31630\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_29\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_30_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31620\,
            in1 => \N__33883\,
            in2 => \_gnd_net_\,
            in3 => \N__31627\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.counter_cry_29\,
            carryout => \phase_controller_inst2.stoper_hc.counter_cry_30\,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst2.stoper_hc.counter_31_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__33898\,
            in1 => \N__31621\,
            in2 => \_gnd_net_\,
            in3 => \N__31495\,
            lcout => \phase_controller_inst2.stoper_hc.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52591\,
            ce => \N__31492\,
            sr => \N__52213\
        );

    \phase_controller_inst1.stoper_tr.counter_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32320\,
            in1 => \N__31426\,
            in2 => \N__31447\,
            in3 => \N__31446\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_0\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32324\,
            in1 => \N__31786\,
            in2 => \_gnd_net_\,
            in3 => \N__31774\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_1\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32321\,
            in1 => \N__31771\,
            in2 => \_gnd_net_\,
            in3 => \N__31759\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_2\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32325\,
            in1 => \N__31756\,
            in2 => \_gnd_net_\,
            in3 => \N__31744\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_3\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32322\,
            in1 => \N__31741\,
            in2 => \_gnd_net_\,
            in3 => \N__31729\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_4\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32326\,
            in1 => \N__31725\,
            in2 => \_gnd_net_\,
            in3 => \N__31711\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_5\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32323\,
            in1 => \N__31708\,
            in2 => \_gnd_net_\,
            in3 => \N__31696\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_6\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_7_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32327\,
            in1 => \N__31692\,
            in2 => \_gnd_net_\,
            in3 => \N__31678\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_7\,
            clk => \N__52586\,
            ce => \N__32191\,
            sr => \N__52220\
        );

    \phase_controller_inst1.stoper_tr.counter_8_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32331\,
            in1 => \N__31675\,
            in2 => \_gnd_net_\,
            in3 => \N__31663\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_8\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_9_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32335\,
            in1 => \N__31660\,
            in2 => \_gnd_net_\,
            in3 => \N__31648\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_9\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_10_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32328\,
            in1 => \N__31932\,
            in2 => \_gnd_net_\,
            in3 => \N__31918\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_10\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_11_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32332\,
            in1 => \N__31915\,
            in2 => \_gnd_net_\,
            in3 => \N__31903\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_11\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_12_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32329\,
            in1 => \N__31900\,
            in2 => \_gnd_net_\,
            in3 => \N__31888\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_12\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_13_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32333\,
            in1 => \N__31885\,
            in2 => \_gnd_net_\,
            in3 => \N__31873\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_13\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_14_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32330\,
            in1 => \N__31870\,
            in2 => \_gnd_net_\,
            in3 => \N__31858\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_14\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_15_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32334\,
            in1 => \N__31855\,
            in2 => \_gnd_net_\,
            in3 => \N__31843\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_15\,
            clk => \N__52581\,
            ce => \N__32190\,
            sr => \N__52229\
        );

    \phase_controller_inst1.stoper_tr.counter_16_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32312\,
            in1 => \N__31827\,
            in2 => \_gnd_net_\,
            in3 => \N__31813\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_16\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_17_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32316\,
            in1 => \N__31803\,
            in2 => \_gnd_net_\,
            in3 => \N__31789\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_17\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_18_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32313\,
            in1 => \N__32066\,
            in2 => \_gnd_net_\,
            in3 => \N__32050\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_18\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_19_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32317\,
            in1 => \N__32045\,
            in2 => \_gnd_net_\,
            in3 => \N__32029\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_19\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_20_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32314\,
            in1 => \N__32096\,
            in2 => \_gnd_net_\,
            in3 => \N__32026\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_20\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_21_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32318\,
            in1 => \N__32114\,
            in2 => \_gnd_net_\,
            in3 => \N__32023\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_21\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_22_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32315\,
            in1 => \N__32708\,
            in2 => \_gnd_net_\,
            in3 => \N__32020\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_22\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_23_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32319\,
            in1 => \N__32741\,
            in2 => \_gnd_net_\,
            in3 => \N__32017\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_23\,
            clk => \N__52576\,
            ce => \N__32189\,
            sr => \N__52235\
        );

    \phase_controller_inst1.stoper_tr.counter_24_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32268\,
            in1 => \N__32007\,
            in2 => \_gnd_net_\,
            in3 => \N__31993\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_24\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_25_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32272\,
            in1 => \N__31983\,
            in2 => \_gnd_net_\,
            in3 => \N__31969\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_25\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_26_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32269\,
            in1 => \N__31953\,
            in2 => \_gnd_net_\,
            in3 => \N__31939\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_26\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_27_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32273\,
            in1 => \N__32361\,
            in2 => \_gnd_net_\,
            in3 => \N__32347\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_27\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_28_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32270\,
            in1 => \N__34543\,
            in2 => \_gnd_net_\,
            in3 => \N__32344\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_28\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_29_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32274\,
            in1 => \N__34558\,
            in2 => \_gnd_net_\,
            in3 => \N__32341\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_29\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_30_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32271\,
            in1 => \N__34504\,
            in2 => \_gnd_net_\,
            in3 => \N__32338\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.counter_cry_29\,
            carryout => \phase_controller_inst1.stoper_tr.counter_cry_30\,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.counter_31_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32275\,
            in1 => \N__34471\,
            in2 => \_gnd_net_\,
            in3 => \N__32194\,
            lcout => \phase_controller_inst1.stoper_tr.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52569\,
            ce => \N__32188\,
            sr => \N__52238\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__32143\,
            in1 => \N__32134\,
            in2 => \N__32122\,
            in3 => \N__32098\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_20_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32161\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52564\,
            ce => \N__36616\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__32142\,
            in1 => \N__32133\,
            in2 => \N__32121\,
            in3 => \N__32097\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__32743\,
            in1 => \N__32725\,
            in2 => \N__32716\,
            in3 => \N__32668\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_22_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32761\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52564\,
            ce => \N__36616\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__32742\,
            in1 => \N__32724\,
            in2 => \N__32715\,
            in3 => \N__32667\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_23_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32686\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52564\,
            ce => \N__36616\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_ticks_28_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34582\,
            lcout => \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52560\,
            ce => \N__32638\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__42556\,
            in1 => \N__51142\,
            in2 => \_gnd_net_\,
            in3 => \N__40039\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32560\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35200\,
            in1 => \N__35363\,
            in2 => \N__35307\,
            in3 => \N__34766\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35857\,
            in1 => \N__35149\,
            in2 => \N__32371\,
            in3 => \N__32938\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32977\,
            in1 => \N__33031\,
            in2 => \N__32965\,
            in3 => \N__32947\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__34946\,
            in1 => \N__34990\,
            in2 => \_gnd_net_\,
            in3 => \N__35041\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__34913\,
            in2 => \N__32956\,
            in3 => \N__32953\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35942\,
            in2 => \_gnd_net_\,
            in3 => \N__35644\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35260\,
            in1 => \N__34823\,
            in2 => \N__32941\,
            in3 => \N__37543\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37696\,
            in1 => \N__37657\,
            in2 => \N__37579\,
            in3 => \N__37609\,
            lcout => \current_shift_inst.PI_CTRL.N_46_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32913\,
            in1 => \N__35866\,
            in2 => \_gnd_net_\,
            in3 => \N__32779\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52551\,
            ce => 'H',
            sr => \N__52248\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35683\,
            in1 => \N__35536\,
            in2 => \N__35616\,
            in3 => \N__35576\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35300\,
            in1 => \N__34759\,
            in2 => \N__35370\,
            in3 => \N__35201\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33022\,
            in1 => \N__33049\,
            in2 => \N__33043\,
            in3 => \N__33016\,
            lcout => \current_shift_inst.PI_CTRL.N_46_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35575\,
            in1 => \N__35611\,
            in2 => \N__35546\,
            in3 => \N__35684\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35472\,
            in1 => \N__35514\,
            in2 => \N__35423\,
            in3 => \N__35893\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34824\,
            in1 => \N__35261\,
            in2 => \N__35953\,
            in3 => \N__35645\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40792\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40633\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40609\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40885\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40813\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40837\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40861\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40909\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52634\,
            ce => \N__41932\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41083\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40744\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41059\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41563\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_18_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40978\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40720\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40768\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52628\,
            ce => \N__41933\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__33280\,
            in1 => \N__33271\,
            in2 => \N__33250\,
            in3 => \N__33214\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_16_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41032\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52622\,
            ce => \N__41934\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__33279\,
            in1 => \N__33270\,
            in2 => \N__33249\,
            in3 => \N__33213\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_17_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41005\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52622\,
            ce => \N__41934\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__33204\,
            in1 => \N__33190\,
            in2 => \N__33165\,
            in3 => \N__33120\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_19_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40956\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52622\,
            ce => \N__41934\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_20_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40930\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52612\,
            ce => \N__41947\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41224\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52612\,
            ce => \N__41947\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_22_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41203\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52612\,
            ce => \N__41947\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_23_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41182\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52612\,
            ce => \N__41947\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__33320\,
            in1 => \N__36147\,
            in2 => \_gnd_net_\,
            in3 => \N__36165\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_28_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42601\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52604\,
            ce => \N__42032\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__33319\,
            in1 => \N__36146\,
            in2 => \_gnd_net_\,
            in3 => \N__36164\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__36104\,
            in1 => \N__36128\,
            in2 => \_gnd_net_\,
            in3 => \N__33321\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__33322\,
            in1 => \N__36105\,
            in2 => \_gnd_net_\,
            in3 => \N__36129\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__33571\,
            in1 => \N__33562\,
            in2 => \N__33543\,
            in3 => \N__33523\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_24_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52597\,
            ce => \N__41948\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__33570\,
            in1 => \N__33561\,
            in2 => \N__33544\,
            in3 => \N__33522\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__33484\,
            in1 => \N__33475\,
            in2 => \N__33457\,
            in3 => \N__33415\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_26_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41122\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52597\,
            ce => \N__41948\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__33483\,
            in1 => \N__33474\,
            in2 => \N__33456\,
            in3 => \N__33414\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_27_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41104\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52597\,
            ce => \N__41948\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__33911\,
            in1 => \N__33393\,
            in2 => \_gnd_net_\,
            in3 => \N__33378\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_28_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42597\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52589\,
            ce => \N__41953\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__33910\,
            in1 => \N__33392\,
            in2 => \_gnd_net_\,
            in3 => \N__33377\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__33896\,
            in1 => \N__33881\,
            in2 => \_gnd_net_\,
            in3 => \N__33912\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__33913\,
            in1 => \N__33897\,
            in2 => \_gnd_net_\,
            in3 => \N__33882\,
            lcout => \phase_controller_inst2.stoper_hc.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47524\,
            in2 => \_gnd_net_\,
            in3 => \N__47501\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__47502\,
            in1 => \_gnd_net_\,
            in2 => \N__47534\,
            in3 => \N__47580\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52585\,
            ce => 'H',
            sr => \N__52208\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__33768\,
            in1 => \N__33850\,
            in2 => \_gnd_net_\,
            in3 => \N__33832\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33826\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33769\,
            in1 => \N__33792\,
            in2 => \_gnd_net_\,
            in3 => \N__33814\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33770\,
            in1 => \N__33592\,
            in2 => \_gnd_net_\,
            in3 => \N__33610\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33586\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_flag_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__34032\,
            in1 => \N__33989\,
            in2 => \N__33973\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52580\,
            ce => 'H',
            sr => \N__52214\
        );

    \phase_controller_inst1.state_4_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__33990\,
            in1 => \N__33968\,
            in2 => \_gnd_net_\,
            in3 => \N__34033\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52580\,
            ce => 'H',
            sr => \N__52214\
        );

    \phase_controller_inst2.start_flag_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__34034\,
            in1 => \_gnd_net_\,
            in2 => \N__34062\,
            in3 => \N__34076\,
            lcout => \phase_controller_inst2.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52580\,
            ce => 'H',
            sr => \N__52214\
        );

    \phase_controller_inst2.state_4_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34077\,
            in1 => \N__34055\,
            in2 => \_gnd_net_\,
            in3 => \N__34035\,
            lcout => \phase_controller_inst2.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52580\,
            ce => 'H',
            sr => \N__52214\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__36409\,
            in1 => \N__50328\,
            in2 => \N__33951\,
            in3 => \N__33933\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.state_ns_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__34036\,
            in1 => \N__33991\,
            in2 => \N__33976\,
            in3 => \N__33972\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52575\,
            ce => 'H',
            sr => \N__52221\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36771\,
            in2 => \_gnd_net_\,
            in3 => \N__36803\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un4_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__34310\,
            in1 => \N__33950\,
            in2 => \N__33955\,
            in3 => \N__34335\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52575\,
            ce => 'H',
            sr => \N__52221\
        );

    \phase_controller_inst1.state_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__36333\,
            in1 => \N__38096\,
            in2 => \N__33952\,
            in3 => \N__33934\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52575\,
            ce => 'H',
            sr => \N__52221\
        );

    \phase_controller_inst1.start_timer_tr_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__38095\,
            in1 => \N__36332\,
            in2 => \N__36780\,
            in3 => \N__36223\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52575\,
            ce => 'H',
            sr => \N__52221\
        );

    \phase_controller_inst1.stoper_tr.running_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__36772\,
            in1 => \N__34311\,
            in2 => \N__36814\,
            in3 => \N__34336\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52575\,
            ce => 'H',
            sr => \N__52221\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34291\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34261\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34234\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34201\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34174\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34141\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34114\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52568\,
            ce => \N__36593\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__34485\,
            in1 => \N__34557\,
            in2 => \_gnd_net_\,
            in3 => \N__34542\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34581\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52562\,
            ce => \N__36595\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__34484\,
            in1 => \N__34556\,
            in2 => \_gnd_net_\,
            in3 => \N__34541\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__34469\,
            in1 => \N__34502\,
            in2 => \_gnd_net_\,
            in3 => \N__34483\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__34503\,
            in1 => \_gnd_net_\,
            in2 => \N__34489\,
            in3 => \N__34470\,
            lcout => \phase_controller_inst1.stoper_tr.un6_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34447\,
            in2 => \_gnd_net_\,
            in3 => \N__34399\,
            lcout => \phase_controller_inst2.stoper_hc.un4_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37404\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52558\,
            ce => 'H',
            sr => \N__52239\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36984\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52558\,
            ce => 'H',
            sr => \N__52239\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37008\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52558\,
            ce => 'H',
            sr => \N__52239\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37233\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52558\,
            ce => 'H',
            sr => \N__52239\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37068\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52554\,
            ce => 'H',
            sr => \N__52241\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37206\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52554\,
            ce => 'H',
            sr => \N__52241\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37179\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52554\,
            ce => 'H',
            sr => \N__52241\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37095\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52554\,
            ce => 'H',
            sr => \N__52241\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37434\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52554\,
            ce => 'H',
            sr => \N__52241\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36957\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52554\,
            ce => 'H',
            sr => \N__52241\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37374\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37041\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37350\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37323\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37296\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37263\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37119\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52549\,
            ce => 'H',
            sr => \N__52243\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34725\,
            in2 => \N__34708\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34675\,
            in2 => \N__34666\,
            in3 => \N__34639\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34636\,
            in2 => \N__34606\,
            in3 => \N__34594\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35110\,
            in2 => \N__35101\,
            in3 => \N__35068\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35065\,
            in2 => \N__35056\,
            in3 => \N__35014\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35011\,
            in2 => \N__35002\,
            in3 => \N__34966\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34963\,
            in2 => \N__34957\,
            in3 => \N__34924\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34921\,
            in2 => \N__34888\,
            in3 => \N__34879\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__52546\,
            ce => 'H',
            sr => \N__52246\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34876\,
            in2 => \N__34867\,
            in3 => \N__34831\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34828\,
            in2 => \N__34798\,
            in3 => \N__34786\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34783\,
            in2 => \N__34774\,
            in3 => \N__34732\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35434\,
            in2 => \N__35425\,
            in3 => \N__35383\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35380\,
            in2 => \N__35371\,
            in3 => \N__35326\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35323\,
            in2 => \N__35314\,
            in3 => \N__35278\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35275\,
            in2 => \N__35266\,
            in3 => \N__35224\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35221\,
            in2 => \N__35212\,
            in3 => \N__35179\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__52543\,
            ce => 'H',
            sr => \N__52249\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35176\,
            in2 => \N__37632\,
            in3 => \N__35167\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37510\,
            in2 => \N__35164\,
            in3 => \N__35128\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35125\,
            in2 => \N__37672\,
            in3 => \N__35113\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37918\,
            in2 => \N__37711\,
            in3 => \N__35698\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37888\,
            in2 => \N__35695\,
            in3 => \N__35665\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37585\,
            in2 => \N__37978\,
            in3 => \N__35662\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37945\,
            in2 => \N__35659\,
            in3 => \N__35626\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37477\,
            in2 => \N__35623\,
            in3 => \N__35590\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__52541\,
            ce => 'H',
            sr => \N__52254\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38188\,
            in2 => \N__35587\,
            in3 => \N__35557\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37771\,
            in2 => \N__35554\,
            in3 => \N__35521\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37801\,
            in2 => \N__35518\,
            in3 => \N__35479\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38161\,
            in2 => \N__35476\,
            in3 => \N__35437\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37828\,
            in2 => \N__35952\,
            in3 => \N__35908\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37861\,
            in2 => \N__35905\,
            in3 => \N__35869\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35862\,
            in1 => \N__38215\,
            in2 => \_gnd_net_\,
            in3 => \N__35722\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52539\,
            ce => 'H',
            sr => \N__52258\
        );

    \GB_BUFFER_reset_c_g_THRU_LUT4_0_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__52294\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_reset_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_16_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41031\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52636\,
            ce => \N__42037\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_17_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41004\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52636\,
            ce => \N__42037\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__35707\,
            in1 => \N__36079\,
            in2 => \N__36057\,
            in3 => \N__35983\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_18_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40977\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52636\,
            ce => \N__42037\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__35706\,
            in1 => \N__36078\,
            in2 => \N__36058\,
            in3 => \N__35982\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_19_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40957\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52636\,
            ce => \N__42037\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.counter_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36922\,
            in1 => \N__38058\,
            in2 => \N__38752\,
            in3 => \N__38751\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_0\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36933\,
            in1 => \N__38031\,
            in2 => \_gnd_net_\,
            in3 => \N__35974\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_1\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36923\,
            in1 => \N__38421\,
            in2 => \_gnd_net_\,
            in3 => \N__35971\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_2\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_3_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36934\,
            in1 => \N__38397\,
            in2 => \_gnd_net_\,
            in3 => \N__35968\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_3\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36924\,
            in1 => \N__38373\,
            in2 => \_gnd_net_\,
            in3 => \N__35965\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_4\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36935\,
            in1 => \N__38349\,
            in2 => \_gnd_net_\,
            in3 => \N__35962\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_5\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36925\,
            in1 => \N__38322\,
            in2 => \_gnd_net_\,
            in3 => \N__35959\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_6\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36936\,
            in1 => \N__38301\,
            in2 => \_gnd_net_\,
            in3 => \N__35956\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_7\,
            clk => \N__52630\,
            ce => \N__36214\,
            sr => \N__52174\
        );

    \phase_controller_inst1.stoper_hc.counter_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36921\,
            in1 => \N__38271\,
            in2 => \_gnd_net_\,
            in3 => \N__36010\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_8\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_9_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36940\,
            in1 => \N__38247\,
            in2 => \_gnd_net_\,
            in3 => \N__36007\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_9\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_10_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36918\,
            in1 => \N__38586\,
            in2 => \_gnd_net_\,
            in3 => \N__36004\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_10\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36937\,
            in1 => \N__38562\,
            in2 => \_gnd_net_\,
            in3 => \N__36001\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_11\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_12_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36919\,
            in1 => \N__38538\,
            in2 => \_gnd_net_\,
            in3 => \N__35998\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_12\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_13_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36938\,
            in1 => \N__38514\,
            in2 => \_gnd_net_\,
            in3 => \N__35995\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_13\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_14_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36920\,
            in1 => \N__38487\,
            in2 => \_gnd_net_\,
            in3 => \N__35992\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_14\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_15_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36939\,
            in1 => \N__38460\,
            in2 => \_gnd_net_\,
            in3 => \N__35989\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_15\,
            clk => \N__52623\,
            ce => \N__36209\,
            sr => \N__52176\
        );

    \phase_controller_inst1.stoper_hc.counter_16_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36914\,
            in1 => \N__38854\,
            in2 => \_gnd_net_\,
            in3 => \N__35986\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_16\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_17_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36929\,
            in1 => \N__38871\,
            in2 => \_gnd_net_\,
            in3 => \N__36082\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_17\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_18_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36915\,
            in1 => \N__36077\,
            in2 => \_gnd_net_\,
            in3 => \N__36061\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_18\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_19_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36930\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__36031\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_19\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_20_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36916\,
            in1 => \N__38720\,
            in2 => \_gnd_net_\,
            in3 => \N__36028\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_20\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_21_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36931\,
            in1 => \N__38737\,
            in2 => \_gnd_net_\,
            in3 => \N__36025\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_21\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_22_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36917\,
            in1 => \N__39023\,
            in2 => \_gnd_net_\,
            in3 => \N__36022\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_22\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_23_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36932\,
            in1 => \N__39049\,
            in2 => \_gnd_net_\,
            in3 => \N__36019\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_23\,
            clk => \N__52615\,
            ce => \N__36213\,
            sr => \N__52179\
        );

    \phase_controller_inst1.stoper_hc.counter_24_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36909\,
            in1 => \N__38951\,
            in2 => \_gnd_net_\,
            in3 => \N__36016\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_24\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_25_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36926\,
            in1 => \N__38968\,
            in2 => \_gnd_net_\,
            in3 => \N__36013\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_25\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_26_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36910\,
            in1 => \N__39112\,
            in2 => \_gnd_net_\,
            in3 => \N__36172\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_26\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_27_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36927\,
            in1 => \N__39136\,
            in2 => \_gnd_net_\,
            in3 => \N__36169\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_27\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_28_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36911\,
            in1 => \N__36166\,
            in2 => \_gnd_net_\,
            in3 => \N__36151\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_28\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_29_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36928\,
            in1 => \N__36148\,
            in2 => \_gnd_net_\,
            in3 => \N__36133\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_29\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_30_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36912\,
            in1 => \N__36130\,
            in2 => \_gnd_net_\,
            in3 => \N__36112\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.counter_cry_29\,
            carryout => \phase_controller_inst1.stoper_hc.counter_cry_30\,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.counter_31_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36106\,
            in1 => \N__36913\,
            in2 => \_gnd_net_\,
            in3 => \N__36109\,
            lcout => \phase_controller_inst1.stoper_hc.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52606\,
            ce => \N__36205\,
            sr => \N__52188\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36249\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50485\,
            in1 => \N__36091\,
            in2 => \_gnd_net_\,
            in3 => \N__46576\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => \elapsed_time_ns_1_RNI36DN9_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36085\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36250\,
            in1 => \_gnd_net_\,
            in2 => \N__50528\,
            in3 => \N__46960\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46927\,
            in1 => \N__36241\,
            in2 => \_gnd_net_\,
            in3 => \N__50484\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36235\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36232\,
            in1 => \N__46996\,
            in2 => \_gnd_net_\,
            in3 => \N__50486\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => \elapsed_time_ns_1_RNI7ADN9_0_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36226\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__36293\,
            in1 => \N__36404\,
            in2 => \N__36274\,
            in3 => \N__50341\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52592\,
            ce => 'H',
            sr => \N__52197\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36292\,
            in2 => \_gnd_net_\,
            in3 => \N__36268\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__36374\,
            in1 => \N__36356\,
            in2 => \_gnd_net_\,
            in3 => \N__38808\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__36358\,
            in1 => \N__36375\,
            in2 => \N__38817\,
            in3 => \N__38775\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52592\,
            ce => 'H',
            sr => \N__52197\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52291\,
            in1 => \N__36357\,
            in2 => \_gnd_net_\,
            in3 => \N__38807\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__36497\,
            in1 => \_gnd_net_\,
            in2 => \N__38155\,
            in3 => \N__38136\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_168_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__38137\,
            in1 => \N__36498\,
            in2 => \_gnd_net_\,
            in3 => \N__38154\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52587\,
            ce => 'H',
            sr => \N__52209\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36496\,
            in2 => \_gnd_net_\,
            in3 => \N__38150\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011001010"
        )
    port map (
            in0 => \N__36354\,
            in1 => \N__50332\,
            in2 => \N__36301\,
            in3 => \N__36405\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52587\,
            ce => 'H',
            sr => \N__52209\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36353\,
            in2 => \_gnd_net_\,
            in3 => \N__38812\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un4_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__36376\,
            in1 => \N__36272\,
            in2 => \N__36361\,
            in3 => \N__38779\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52587\,
            ce => 'H',
            sr => \N__52209\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36355\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52587\,
            ce => 'H',
            sr => \N__52209\
        );

    \phase_controller_inst1.state_1_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__36334\,
            in1 => \N__36300\,
            in2 => \N__38100\,
            in3 => \N__36273\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52582\,
            ce => 'H',
            sr => \N__52215\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36776\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52582\,
            ce => 'H',
            sr => \N__52215\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38816\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__36802\,
            in1 => \N__52293\,
            in2 => \_gnd_net_\,
            in3 => \N__36770\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48116\,
            in1 => \N__49494\,
            in2 => \N__50113\,
            in3 => \N__48097\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48115\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47887\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47758\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_ticks_0_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36741\,
            in2 => \_gnd_net_\,
            in3 => \N__36703\,
            lcout => \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52570\,
            ce => \N__36594\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47275\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44669\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44044\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44561\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48050\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47986\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44443\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37024\,
            in2 => \_gnd_net_\,
            in3 => \N__40030\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40021\,
            in2 => \_gnd_net_\,
            in3 => \N__36994\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40009\,
            in2 => \_gnd_net_\,
            in3 => \N__36970\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39997\,
            in2 => \_gnd_net_\,
            in3 => \N__36943\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39985\,
            in2 => \_gnd_net_\,
            in3 => \N__37219\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39970\,
            in2 => \_gnd_net_\,
            in3 => \N__37192\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40153\,
            in3 => \N__37165\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40138\,
            in2 => \_gnd_net_\,
            in3 => \N__37132\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__52565\,
            ce => 'H',
            sr => \N__52236\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40126\,
            in2 => \_gnd_net_\,
            in3 => \N__37105\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40114\,
            in2 => \_gnd_net_\,
            in3 => \N__37081\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40102\,
            in2 => \_gnd_net_\,
            in3 => \N__37054\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40090\,
            in2 => \_gnd_net_\,
            in3 => \N__37027\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40078\,
            in2 => \_gnd_net_\,
            in3 => \N__37420\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40066\,
            in2 => \_gnd_net_\,
            in3 => \N__37390\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40054\,
            in3 => \N__37360\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40252\,
            in2 => \_gnd_net_\,
            in3 => \N__37336\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__52561\,
            ce => 'H',
            sr => \N__52240\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40240\,
            in2 => \_gnd_net_\,
            in3 => \N__37309\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40228\,
            in2 => \_gnd_net_\,
            in3 => \N__37282\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40216\,
            in2 => \_gnd_net_\,
            in3 => \N__37279\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40204\,
            in2 => \_gnd_net_\,
            in3 => \N__37249\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40192\,
            in2 => \_gnd_net_\,
            in3 => \N__37246\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40180\,
            in2 => \_gnd_net_\,
            in3 => \N__37471\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40168\,
            in3 => \N__37468\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40348\,
            in2 => \_gnd_net_\,
            in3 => \N__37465\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__52556\,
            ce => 'H',
            sr => \N__52242\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40336\,
            in2 => \_gnd_net_\,
            in3 => \N__37462\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40324\,
            in2 => \_gnd_net_\,
            in3 => \N__37459\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40312\,
            in2 => \_gnd_net_\,
            in3 => \N__37456\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40300\,
            in2 => \_gnd_net_\,
            in3 => \N__37453\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40288\,
            in2 => \_gnd_net_\,
            in3 => \N__37450\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40276\,
            in2 => \_gnd_net_\,
            in3 => \N__37447\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40522\,
            in3 => \N__37765\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40261\,
            in2 => \_gnd_net_\,
            in3 => \N__37762\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52552\,
            ce => 'H',
            sr => \N__52244\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37750\,
            in1 => \N__37759\,
            in2 => \N__37732\,
            in3 => \N__37740\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37758\,
            in1 => \N__40440\,
            in2 => \N__40468\,
            in3 => \N__37749\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40503\,
            in2 => \_gnd_net_\,
            in3 => \N__40482\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37741\,
            in1 => \N__37731\,
            in2 => \N__37720\,
            in3 => \N__37717\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37703\,
            in1 => \N__37671\,
            in2 => \N__37633\,
            in3 => \N__37584\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52544\,
            ce => 'H',
            sr => \N__52250\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37497\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52544\,
            ce => 'H',
            sr => \N__52250\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38004\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52544\,
            ce => 'H',
            sr => \N__52250\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37962\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52544\,
            ce => 'H',
            sr => \N__52250\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37938\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52544\,
            ce => 'H',
            sr => \N__52250\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37908\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52544\,
            ce => 'H',
            sr => \N__52250\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37878\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37848\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37821\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37788\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38224\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38205\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38181\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52542\,
            ce => 'H',
            sr => \N__52255\
        );

    \delay_measurement_inst.stop_timer_tr_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38127\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38110\,
            ce => 'H',
            sr => \N__52259\
        );

    \delay_measurement_inst.start_timer_tr_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38126\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38110\,
            ce => 'H',
            sr => \N__52259\
        );

    \phase_controller_inst1.S2_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38101\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52538\,
            ce => 'H',
            sr => \N__52265\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40696\,
            in2 => \N__38044\,
            in3 => \N__38062\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40555\,
            in2 => \N__38017\,
            in3 => \N__38035\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38407\,
            in2 => \N__40357\,
            in3 => \N__38422\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38401\,
            in1 => \N__40576\,
            in2 => \N__38383\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38359\,
            in2 => \N__40564\,
            in3 => \N__38374\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40549\,
            in2 => \N__38335\,
            in3 => \N__38353\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38308\,
            in2 => \N__40585\,
            in3 => \N__38326\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38302\,
            in1 => \N__40570\,
            in2 => \N__38287\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40669\,
            in2 => \N__38257\,
            in3 => \N__38275\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40675\,
            in2 => \N__38233\,
            in3 => \N__38248\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40681\,
            in2 => \N__38572\,
            in3 => \N__38590\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40537\,
            in2 => \N__38548\,
            in3 => \N__38563\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38524\,
            in2 => \N__40690\,
            in3 => \N__38539\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40543\,
            in2 => \N__38500\,
            in3 => \N__38518\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38488\,
            in1 => \N__40531\,
            in2 => \N__38473\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38464\,
            in1 => \N__41542\,
            in2 => \N__38446\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.counter_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38596\,
            in2 => \N__38839\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38437\,
            in2 => \N__38431\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38602\,
            in2 => \N__38701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39004\,
            in2 => \N__38674\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38986\,
            in2 => \N__38932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38911\,
            in2 => \N__39097\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38662\,
            in2 => \N__38650\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38635\,
            in2 => \N__38620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un6_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un6_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38605\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__38691\,
            in1 => \N__38735\,
            in2 => \N__38721\,
            in3 => \N__38682\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__38853\,
            in1 => \N__38870\,
            in2 => \N__38887\,
            in3 => \N__38902\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__38901\,
            in1 => \N__38886\,
            in2 => \N__38872\,
            in3 => \N__38852\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43711\,
            in1 => \N__50529\,
            in2 => \_gnd_net_\,
            in3 => \N__38827\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => \elapsed_time_ns_1_RNIG23T9_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38821\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38818\,
            in2 => \_gnd_net_\,
            in3 => \N__38763\,
            lcout => \phase_controller_inst1.stoper_hc.counter\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__38692\,
            in1 => \N__38736\,
            in2 => \N__38722\,
            in3 => \N__38683\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_20_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40923\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52624\,
            ce => \N__42033\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_21_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41217\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52624\,
            ce => \N__42033\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__39048\,
            in1 => \N__39034\,
            in2 => \N__39025\,
            in3 => \N__38995\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_22_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41196\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52624\,
            ce => \N__42033\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__39047\,
            in1 => \N__39033\,
            in2 => \N__39024\,
            in3 => \N__38994\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_23_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41175\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52624\,
            ce => \N__42033\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__38977\,
            in1 => \N__38967\,
            in2 => \N__38953\,
            in3 => \N__38920\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_24_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41157\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52616\,
            ce => \N__42022\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__38976\,
            in1 => \N__38966\,
            in2 => \N__38952\,
            in3 => \N__38919\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_25_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41136\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52616\,
            ce => \N__42022\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__39135\,
            in1 => \N__39121\,
            in2 => \N__39085\,
            in3 => \N__39111\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_26_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41118\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52616\,
            ce => \N__42022\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__39134\,
            in1 => \N__39120\,
            in2 => \N__39084\,
            in3 => \N__39110\,
            lcout => \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_27_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41100\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52616\,
            ce => \N__42022\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47246\,
            in1 => \N__42521\,
            in2 => \_gnd_net_\,
            in3 => \N__39070\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_1_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47238\,
            in1 => \N__41243\,
            in2 => \_gnd_net_\,
            in3 => \N__39067\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_2_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47247\,
            in1 => \N__39237\,
            in2 => \_gnd_net_\,
            in3 => \N__39064\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_3_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47239\,
            in1 => \N__39209\,
            in2 => \_gnd_net_\,
            in3 => \N__39061\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_4_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47248\,
            in1 => \N__39507\,
            in2 => \_gnd_net_\,
            in3 => \N__39058\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_5_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47240\,
            in1 => \N__39482\,
            in2 => \_gnd_net_\,
            in3 => \N__39055\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_6_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47249\,
            in1 => \N__39450\,
            in2 => \_gnd_net_\,
            in3 => \N__39052\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_7_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47241\,
            in1 => \N__39422\,
            in2 => \_gnd_net_\,
            in3 => \N__39163\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__52607\,
            ce => \N__47367\,
            sr => \N__52189\
        );

    \current_shift_inst.timer_s1.counter_8_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47237\,
            in1 => \N__39398\,
            in2 => \_gnd_net_\,
            in3 => \N__39160\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_9_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47245\,
            in1 => \N__39368\,
            in2 => \_gnd_net_\,
            in3 => \N__39157\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_10_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47234\,
            in1 => \N__39335\,
            in2 => \_gnd_net_\,
            in3 => \N__39154\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_11_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47242\,
            in1 => \N__39309\,
            in2 => \_gnd_net_\,
            in3 => \N__39151\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_12_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47235\,
            in1 => \N__39285\,
            in2 => \_gnd_net_\,
            in3 => \N__39148\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_13_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47243\,
            in1 => \N__39719\,
            in2 => \_gnd_net_\,
            in3 => \N__39145\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_14_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47236\,
            in1 => \N__39687\,
            in2 => \_gnd_net_\,
            in3 => \N__39142\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_15_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47244\,
            in1 => \N__39665\,
            in2 => \_gnd_net_\,
            in3 => \N__39139\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__52599\,
            ce => \N__47360\,
            sr => \N__52192\
        );

    \current_shift_inst.timer_s1.counter_16_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47254\,
            in1 => \N__39635\,
            in2 => \_gnd_net_\,
            in3 => \N__39190\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_17_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47250\,
            in1 => \N__39605\,
            in2 => \_gnd_net_\,
            in3 => \N__39187\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_18_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47255\,
            in1 => \N__39581\,
            in2 => \_gnd_net_\,
            in3 => \N__39184\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_19_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47251\,
            in1 => \N__39560\,
            in2 => \_gnd_net_\,
            in3 => \N__39181\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_20_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47256\,
            in1 => \N__39533\,
            in2 => \_gnd_net_\,
            in3 => \N__39178\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_21_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47252\,
            in1 => \N__39950\,
            in2 => \_gnd_net_\,
            in3 => \N__39175\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_22_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47257\,
            in1 => \N__39924\,
            in2 => \_gnd_net_\,
            in3 => \N__39172\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_23_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47253\,
            in1 => \N__39896\,
            in2 => \_gnd_net_\,
            in3 => \N__39169\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__52593\,
            ce => \N__47371\,
            sr => \N__52198\
        );

    \current_shift_inst.timer_s1.counter_24_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47228\,
            in1 => \N__39869\,
            in2 => \_gnd_net_\,
            in3 => \N__39166\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__52588\,
            ce => \N__47353\,
            sr => \N__52210\
        );

    \current_shift_inst.timer_s1.counter_25_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47232\,
            in1 => \N__39839\,
            in2 => \_gnd_net_\,
            in3 => \N__39268\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__52588\,
            ce => \N__47353\,
            sr => \N__52210\
        );

    \current_shift_inst.timer_s1.counter_26_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47229\,
            in1 => \N__39797\,
            in2 => \_gnd_net_\,
            in3 => \N__39265\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__52588\,
            ce => \N__47353\,
            sr => \N__52210\
        );

    \current_shift_inst.timer_s1.counter_27_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47233\,
            in1 => \N__39752\,
            in2 => \_gnd_net_\,
            in3 => \N__39262\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__52588\,
            ce => \N__47353\,
            sr => \N__52210\
        );

    \current_shift_inst.timer_s1.counter_28_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47230\,
            in1 => \N__39816\,
            in2 => \_gnd_net_\,
            in3 => \N__39259\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__52588\,
            ce => \N__47353\,
            sr => \N__52210\
        );

    \current_shift_inst.timer_s1.counter_29_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__39771\,
            in1 => \N__47231\,
            in2 => \_gnd_net_\,
            in3 => \N__39256\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52588\,
            ce => \N__47353\,
            sr => \N__52210\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42525\,
            in2 => \N__39249\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41245\,
            in2 => \N__39220\,
            in3 => \N__39253\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39513\,
            in2 => \N__39250\,
            in3 => \N__39223\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39219\,
            in2 => \N__39489\,
            in3 => \N__39193\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39514\,
            in2 => \N__39462\,
            in3 => \N__39493\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39429\,
            in2 => \N__39490\,
            in3 => \N__39466\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39399\,
            in2 => \N__39463\,
            in3 => \N__39436\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39369\,
            in2 => \N__39433\,
            in3 => \N__39406\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__52583\,
            ce => \N__44194\,
            sr => \N__52216\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39342\,
            in2 => \N__39403\,
            in3 => \N__39379\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39315\,
            in2 => \N__39376\,
            in3 => \N__39349\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39291\,
            in2 => \N__39346\,
            in3 => \N__39319\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39316\,
            in2 => \N__39726\,
            in3 => \N__39295\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39292\,
            in2 => \N__39699\,
            in3 => \N__39271\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39666\,
            in2 => \N__39727\,
            in3 => \N__39703\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39636\,
            in2 => \N__39700\,
            in3 => \N__39673\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39606\,
            in2 => \N__39670\,
            in3 => \N__39646\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__52577\,
            ce => \N__44193\,
            sr => \N__52222\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39582\,
            in2 => \N__39643\,
            in3 => \N__39616\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39561\,
            in2 => \N__39613\,
            in3 => \N__39586\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39583\,
            in2 => \N__39540\,
            in3 => \N__39565\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39562\,
            in2 => \N__39957\,
            in3 => \N__39544\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39930\,
            in2 => \N__39541\,
            in3 => \N__39517\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39903\,
            in2 => \N__39958\,
            in3 => \N__39934\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39931\,
            in2 => \N__39876\,
            in3 => \N__39910\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39840\,
            in2 => \N__39907\,
            in3 => \N__39880\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__52571\,
            ce => \N__44192\,
            sr => \N__52230\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39798\,
            in2 => \N__39877\,
            in3 => \N__39850\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__52566\,
            ce => \N__44191\,
            sr => \N__52237\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39753\,
            in2 => \N__39847\,
            in3 => \N__39820\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__52566\,
            ce => \N__44191\,
            sr => \N__52237\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39817\,
            in2 => \N__39802\,
            in3 => \N__39778\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__52566\,
            ce => \N__44191\,
            sr => \N__52237\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39775\,
            in2 => \N__39757\,
            in3 => \N__39733\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__52566\,
            ce => \N__44191\,
            sr => \N__52237\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39730\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44371\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43396\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44213\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52566\,
            ce => \N__44191\,
            sr => \N__52237\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43102\,
            in2 => \N__43090\,
            in3 => \N__43089\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41461\,
            in2 => \_gnd_net_\,
            in3 => \N__40012\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41455\,
            in2 => \_gnd_net_\,
            in3 => \N__40000\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41449\,
            in2 => \_gnd_net_\,
            in3 => \N__39988\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41443\,
            in2 => \_gnd_net_\,
            in3 => \N__39973\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41437\,
            in2 => \_gnd_net_\,
            in3 => \N__39961\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41431\,
            in2 => \_gnd_net_\,
            in3 => \N__40141\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41533\,
            in2 => \_gnd_net_\,
            in3 => \N__40129\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43300\,
            in2 => \_gnd_net_\,
            in3 => \N__40117\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43114\,
            in2 => \_gnd_net_\,
            in3 => \N__40105\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43066\,
            in2 => \_gnd_net_\,
            in3 => \N__40093\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43312\,
            in2 => \_gnd_net_\,
            in3 => \N__40081\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43273\,
            in2 => \_gnd_net_\,
            in3 => \N__40069\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41527\,
            in2 => \_gnd_net_\,
            in3 => \N__40057\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43291\,
            in2 => \_gnd_net_\,
            in3 => \N__40042\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43282\,
            in2 => \_gnd_net_\,
            in3 => \N__40243\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41497\,
            in2 => \_gnd_net_\,
            in3 => \N__40231\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41503\,
            in2 => \_gnd_net_\,
            in3 => \N__40219\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41668\,
            in2 => \_gnd_net_\,
            in3 => \N__40207\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43510\,
            in2 => \_gnd_net_\,
            in3 => \N__40195\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43429\,
            in2 => \_gnd_net_\,
            in3 => \N__40183\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41521\,
            in2 => \_gnd_net_\,
            in3 => \N__40171\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41509\,
            in2 => \_gnd_net_\,
            in3 => \N__40156\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49039\,
            in2 => \_gnd_net_\,
            in3 => \N__40339\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43264\,
            in2 => \_gnd_net_\,
            in3 => \N__40327\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41491\,
            in2 => \_gnd_net_\,
            in3 => \N__40315\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41515\,
            in2 => \_gnd_net_\,
            in3 => \N__40303\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41485\,
            in2 => \_gnd_net_\,
            in3 => \N__40291\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45367\,
            in2 => \_gnd_net_\,
            in3 => \N__40279\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41767\,
            in2 => \_gnd_net_\,
            in3 => \N__40267\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49164\,
            in2 => \_gnd_net_\,
            in3 => \N__40264\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => \current_shift_inst.control_input_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40525\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41646\,
            in2 => \_gnd_net_\,
            in3 => \N__41625\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40392\,
            in1 => \N__40377\,
            in2 => \N__40510\,
            in3 => \N__40407\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41761\,
            in1 => \N__40507\,
            in2 => \N__40489\,
            in3 => \N__41740\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40422\,
            in1 => \N__40467\,
            in2 => \N__40447\,
            in3 => \N__41661\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40426\,
            in1 => \N__40408\,
            in2 => \N__40396\,
            in3 => \N__40378\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47563\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40366\,
            ce => 'H',
            sr => \N__52168\
        );

    \delay_measurement_inst.stop_timer_hc_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47564\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40366\,
            ce => 'H',
            sr => \N__52168\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40629\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40857\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_3_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40605\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_7_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40833\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_4_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40905\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40653\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_5_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40881\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52653\,
            ce => \N__42043\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_13_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41079\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40740\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_14_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41055\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_0_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42640\,
            in2 => \_gnd_net_\,
            in3 => \N__41833\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40716\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_10_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40764\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_9_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40788\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40812\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52647\,
            ce => \N__42039\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42631\,
            in1 => \N__40663\,
            in2 => \N__41832\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__41796\,
            in2 => \N__51646\,
            in3 => \N__40636\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_1,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41782\,
            in1 => \N__41781\,
            in2 => \N__51659\,
            in3 => \N__40612\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_2,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42175\,
            in1 => \N__42174\,
            in2 => \N__51647\,
            in3 => \N__40588\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_3,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42160\,
            in1 => \N__42159\,
            in2 => \N__51660\,
            in3 => \N__40888\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_4,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42145\,
            in1 => \N__42144\,
            in2 => \N__51648\,
            in3 => \N__40864\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_5,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42130\,
            in1 => \N__42129\,
            in2 => \N__51661\,
            in3 => \N__40840\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_6,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42109\,
            in1 => \N__42108\,
            in2 => \N__51649\,
            in3 => \N__40816\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_7,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42088\,
            in1 => \N__42087\,
            in2 => \N__51590\,
            in3 => \N__40795\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_8,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42073\,
            in1 => \N__42072\,
            in2 => \N__51587\,
            in3 => \N__40771\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_9,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42058\,
            in1 => \N__42057\,
            in2 => \N__51591\,
            in3 => \N__40747\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_10,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42340\,
            in1 => \N__42339\,
            in2 => \N__51584\,
            in3 => \N__40723\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_11,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42325\,
            in1 => \N__42324\,
            in2 => \N__51588\,
            in3 => \N__40699\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_12,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42310\,
            in1 => \N__42309\,
            in2 => \N__51585\,
            in3 => \N__41062\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_13,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42295\,
            in1 => \N__42294\,
            in2 => \N__51589\,
            in3 => \N__41038\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_14,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42274\,
            in1 => \N__42273\,
            in2 => \N__51586\,
            in3 => \N__41035\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_15,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42256\,
            in1 => \N__42255\,
            in2 => \N__51580\,
            in3 => \N__41008\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_16,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42241\,
            in1 => \N__42240\,
            in2 => \N__51604\,
            in3 => \N__40981\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_17,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42219\,
            in1 => \N__42226\,
            in2 => \N__51581\,
            in3 => \N__40960\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_18,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42190\,
            in1 => \N__42189\,
            in2 => \N__51605\,
            in3 => \N__40933\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_19,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42502\,
            in1 => \N__42498\,
            in2 => \N__51582\,
            in3 => \N__40912\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_20,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42484\,
            in1 => \N__42483\,
            in2 => \N__51606\,
            in3 => \N__41206\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_21,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42460\,
            in1 => \N__42459\,
            in2 => \N__51583\,
            in3 => \N__41185\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_22,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42439\,
            in1 => \N__42438\,
            in2 => \N__51607\,
            in3 => \N__41164\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_23,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42421\,
            in1 => \N__42420\,
            in2 => \N__51418\,
            in3 => \N__41146\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_24,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42406\,
            in1 => \N__42405\,
            in2 => \N__51420\,
            in3 => \N__41125\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_25,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42382\,
            in1 => \N__42381\,
            in2 => \N__51419\,
            in3 => \N__41107\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_26,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42355\,
            in1 => \N__42354\,
            in2 => \N__51421\,
            in3 => \N__41089\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_27,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41086\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41256\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43725\,
            in1 => \N__41268\,
            in2 => \N__43710\,
            in3 => \N__46659\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__43849\,
            in1 => \N__41275\,
            in2 => \N__43825\,
            in3 => \N__42580\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45319\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52617\,
            ce => \N__43959\,
            sr => \N__52180\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45685\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52617\,
            ce => \N__43959\,
            sr => \N__52180\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41862\,
            in1 => \N__41269\,
            in2 => \_gnd_net_\,
            in3 => \N__50479\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50480\,
            in1 => \N__41257\,
            in2 => \_gnd_net_\,
            in3 => \N__43729\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__49446\,
            in1 => \N__48327\,
            in2 => \N__48223\,
            in3 => \N__48303\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41244\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52608\,
            ce => \N__44196\,
            sr => \N__52190\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48301\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__43177\,
            in1 => \N__48326\,
            in2 => \_gnd_net_\,
            in3 => \N__48302\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49447\,
            in2 => \_gnd_net_\,
            in3 => \N__44706\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__50754\,
            in1 => \N__49448\,
            in2 => \N__50112\,
            in3 => \N__44707\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44149\,
            in1 => \N__43178\,
            in2 => \_gnd_net_\,
            in3 => \N__44160\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44513\,
            in1 => \N__43182\,
            in2 => \_gnd_net_\,
            in3 => \N__44477\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43183\,
            in1 => \N__47633\,
            in2 => \_gnd_net_\,
            in3 => \N__47660\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48243\,
            in1 => \N__43184\,
            in2 => \_gnd_net_\,
            in3 => \N__48264\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43181\,
            in1 => \N__48386\,
            in2 => \_gnd_net_\,
            in3 => \N__48350\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43179\,
            in1 => \N__46794\,
            in2 => \_gnd_net_\,
            in3 => \N__46764\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__47315\,
            in1 => \N__43180\,
            in2 => \_gnd_net_\,
            in3 => \N__47285\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48242\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44265\,
            in1 => \N__43219\,
            in2 => \_gnd_net_\,
            in3 => \N__44243\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43220\,
            in1 => \N__47063\,
            in2 => \_gnd_net_\,
            in3 => \N__47037\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44503\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46787\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48117\,
            in1 => \N__43218\,
            in2 => \_gnd_net_\,
            in3 => \N__48083\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44135\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47623\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__48372\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44045\,
            in1 => \N__43221\,
            in2 => \_gnd_net_\,
            in3 => \N__44021\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43222\,
            in1 => \N__47720\,
            in2 => \_gnd_net_\,
            in3 => \N__47687\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47412\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47054\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47088\,
            in1 => \N__43223\,
            in2 => \_gnd_net_\,
            in3 => \N__47123\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47087\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47719\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44264\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50744\,
            in2 => \N__42555\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51405\,
            in2 => \N__41296\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41284\,
            in2 => \N__51502\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51409\,
            in2 => \N__41383\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41371\,
            in2 => \N__51503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51413\,
            in2 => \N__41362\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41350\,
            in2 => \N__51504\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51417\,
            in2 => \N__41341\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51401\,
            in2 => \N__41329\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41317\,
            in2 => \N__51501\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51389\,
            in2 => \N__41308\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41425\,
            in2 => \N__51498\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51393\,
            in2 => \N__41416\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41404\,
            in2 => \N__51499\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51397\,
            in2 => \N__41395\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42931\,
            in2 => \N__51500\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51338\,
            in2 => \N__43027\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51342\,
            in2 => \N__42925\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51339\,
            in2 => \N__42574\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51343\,
            in2 => \N__43018\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51340\,
            in2 => \N__42913\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51344\,
            in2 => \N__43036\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51341\,
            in2 => \N__43054\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51345\,
            in2 => \N__43003\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51220\,
            in2 => \N__43126\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43045\,
            in2 => \N__51386\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51224\,
            in2 => \N__42994\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43252\,
            in2 => \N__51387\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51228\,
            in2 => \N__42985\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42976\,
            in2 => \N__51388\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51232\,
            in2 => \N__41479\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49496\,
            in2 => \_gnd_net_\,
            in3 => \N__41464\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48136\,
            in1 => \N__44944\,
            in2 => \_gnd_net_\,
            in3 => \N__49109\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__49110\,
            in1 => \N__48577\,
            in2 => \_gnd_net_\,
            in3 => \N__44917\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48553\,
            in1 => \N__44902\,
            in2 => \_gnd_net_\,
            in3 => \N__49111\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__49112\,
            in1 => \N__44887\,
            in2 => \_gnd_net_\,
            in3 => \N__48529\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__44857\,
            in1 => \N__48499\,
            in2 => \_gnd_net_\,
            in3 => \N__49113\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__49114\,
            in1 => \N__44833\,
            in2 => \_gnd_net_\,
            in3 => \N__48472\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48445\,
            in1 => \N__44803\,
            in2 => \_gnd_net_\,
            in3 => \N__49115\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__49116\,
            in1 => \N__45034\,
            in2 => \_gnd_net_\,
            in3 => \N__48685\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__45178\,
            in1 => \N__48865\,
            in2 => \_gnd_net_\,
            in3 => \N__49157\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__49160\,
            in1 => \N__50155\,
            in2 => \_gnd_net_\,
            in3 => \N__45430\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__45160\,
            in1 => \N__48841\,
            in2 => \_gnd_net_\,
            in3 => \N__49158\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__49156\,
            in1 => \N__48970\,
            in2 => \_gnd_net_\,
            in3 => \N__45277\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__44968\,
            in1 => \N__48604\,
            in2 => \_gnd_net_\,
            in3 => \N__49155\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__49159\,
            in1 => \N__50179\,
            in2 => \_gnd_net_\,
            in3 => \N__45451\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__49161\,
            in1 => \N__50128\,
            in2 => \_gnd_net_\,
            in3 => \N__45397\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41688\,
            in2 => \_gnd_net_\,
            in3 => \N__41760\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41716\,
            in1 => \N__41739\,
            in2 => \N__41719\,
            in3 => \N__41704\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41715\,
            in2 => \_gnd_net_\,
            in3 => \N__41703\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41689\,
            in1 => \N__41607\,
            in2 => \N__41677\,
            in3 => \N__41674\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__45250\,
            in1 => \N__48943\,
            in2 => \_gnd_net_\,
            in3 => \N__49162\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41662\,
            in1 => \N__41647\,
            in2 => \N__41632\,
            in3 => \N__41611\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41590\,
            in1 => \N__41584\,
            in2 => \N__41572\,
            in3 => \N__41569\,
            lcout => \current_shift_inst.PI_CTRL.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41559\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52654\,
            ce => \N__42038\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46702\,
            in1 => \N__42635\,
            in2 => \_gnd_net_\,
            in3 => \N__50547\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => \elapsed_time_ns_1_RNI04EN9_0_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_ticks_0_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41968\,
            in3 => \N__41831\,
            lcout => \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52648\,
            ce => \N__41952\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43579\,
            in1 => \N__46978\,
            in2 => \_gnd_net_\,
            in3 => \N__50548\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42630\,
            in2 => \N__41875\,
            in3 => \N__46648\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41848\,
            in2 => \_gnd_net_\,
            in3 => \N__41866\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41842\,
            in2 => \_gnd_net_\,
            in3 => \N__41809\,
            lcout => \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41806\,
            in2 => \_gnd_net_\,
            in3 => \N__41785\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43516\,
            in2 => \_gnd_net_\,
            in3 => \N__41770\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43774\,
            in2 => \_gnd_net_\,
            in3 => \N__42163\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43588\,
            in2 => \_gnd_net_\,
            in3 => \N__42148\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43663\,
            in2 => \_gnd_net_\,
            in3 => \N__42133\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43633\,
            in2 => \_gnd_net_\,
            in3 => \N__42112\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43678\,
            in2 => \_gnd_net_\,
            in3 => \N__42091\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43759\,
            in2 => \_gnd_net_\,
            in3 => \N__42076\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43627\,
            in2 => \_gnd_net_\,
            in3 => \N__42061\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49003\,
            in2 => \_gnd_net_\,
            in3 => \N__42046\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48994\,
            in2 => \_gnd_net_\,
            in3 => \N__42328\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43744\,
            in2 => \_gnd_net_\,
            in3 => \N__42313\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43648\,
            in2 => \_gnd_net_\,
            in3 => \N__42298\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43555\,
            in2 => \_gnd_net_\,
            in3 => \N__42277\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46537\,
            in2 => \_gnd_net_\,
            in3 => \N__42259\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46717\,
            in2 => \_gnd_net_\,
            in3 => \N__42244\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43534\,
            in2 => \_gnd_net_\,
            in3 => \N__42229\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47593\,
            in2 => \_gnd_net_\,
            in3 => \N__42205\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42202\,
            in2 => \_gnd_net_\,
            in3 => \N__42178\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50629\,
            in2 => \_gnd_net_\,
            in3 => \N__42487\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43567\,
            in2 => \_gnd_net_\,
            in3 => \N__42472\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42469\,
            in2 => \_gnd_net_\,
            in3 => \N__42442\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50605\,
            in2 => \_gnd_net_\,
            in3 => \N__42424\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45346\,
            in2 => \_gnd_net_\,
            in3 => \N__42409\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46237\,
            in2 => \_gnd_net_\,
            in3 => \N__42394\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42391\,
            in2 => \_gnd_net_\,
            in3 => \N__42370\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42367\,
            in2 => \_gnd_net_\,
            in3 => \N__42343\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29\,
            carryout => \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__42646\,
            in1 => \N__42639\,
            in2 => \_gnd_net_\,
            in3 => \N__42604\,
            lcout => phase_controller_inst1_stoper_hc_target_ticks_1_i_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__43878\,
            in1 => \N__43863\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__49497\,
            in1 => \N__47869\,
            in2 => \N__47830\,
            in3 => \N__50077\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__49498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50076\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47868\,
            in1 => \N__43176\,
            in2 => \_gnd_net_\,
            in3 => \N__47825\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44077\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__44078\,
            in1 => \_gnd_net_\,
            in2 => \N__42559\,
            in3 => \N__43175\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44230\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52618\,
            ce => \N__44197\,
            sr => \N__52181\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42529\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52618\,
            ce => \N__44197\,
            sr => \N__52181\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42721\,
            in2 => \N__44118\,
            in3 => \N__44114\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42715\,
            in2 => \_gnd_net_\,
            in3 => \N__42709\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42706\,
            in2 => \_gnd_net_\,
            in3 => \N__42700\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42697\,
            in2 => \_gnd_net_\,
            in3 => \N__42691\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42688\,
            in2 => \_gnd_net_\,
            in3 => \N__42682\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42679\,
            in2 => \_gnd_net_\,
            in3 => \N__42673\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42670\,
            in2 => \_gnd_net_\,
            in3 => \N__42664\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42661\,
            in2 => \_gnd_net_\,
            in3 => \N__42649\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42823\,
            in2 => \_gnd_net_\,
            in3 => \N__42817\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42814\,
            in2 => \_gnd_net_\,
            in3 => \N__42808\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42805\,
            in2 => \_gnd_net_\,
            in3 => \N__42793\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42790\,
            in2 => \_gnd_net_\,
            in3 => \N__42778\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42775\,
            in2 => \_gnd_net_\,
            in3 => \N__42769\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42766\,
            in2 => \_gnd_net_\,
            in3 => \N__42760\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42757\,
            in2 => \_gnd_net_\,
            in3 => \N__42745\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42742\,
            in2 => \_gnd_net_\,
            in3 => \N__42736\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42733\,
            in2 => \_gnd_net_\,
            in3 => \N__42724\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44005\,
            in2 => \_gnd_net_\,
            in3 => \N__42904\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42901\,
            in2 => \_gnd_net_\,
            in3 => \N__42892\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42889\,
            in2 => \_gnd_net_\,
            in3 => \N__42877\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42874\,
            in2 => \_gnd_net_\,
            in3 => \N__42862\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42859\,
            in2 => \_gnd_net_\,
            in3 => \N__42847\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42844\,
            in2 => \_gnd_net_\,
            in3 => \N__42832\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46816\,
            in2 => \_gnd_net_\,
            in3 => \N__42829\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43009\,
            in2 => \_gnd_net_\,
            in3 => \N__42826\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43438\,
            in2 => \_gnd_net_\,
            in3 => \N__42970\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42967\,
            in2 => \_gnd_net_\,
            in3 => \N__42955\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42952\,
            in2 => \_gnd_net_\,
            in3 => \N__42940\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43246\,
            in2 => \_gnd_net_\,
            in3 => \N__42937\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42934\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43229\,
            in1 => \N__44453\,
            in2 => \_gnd_net_\,
            in3 => \N__44414\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__47897\,
            in1 => \N__47930\,
            in2 => \_gnd_net_\,
            in3 => \N__43230\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__49877\,
            in1 => \N__49453\,
            in2 => \N__44526\,
            in3 => \N__44485\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43233\,
            in1 => \N__44676\,
            in2 => \_gnd_net_\,
            in3 => \N__44654\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48059\,
            in1 => \N__43235\,
            in2 => \_gnd_net_\,
            in3 => \N__48033\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__49452\,
            in1 => \N__44723\,
            in2 => \_gnd_net_\,
            in3 => \N__44766\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44568\,
            in1 => \N__43234\,
            in2 => \_gnd_net_\,
            in3 => \N__44547\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__43231\,
            in1 => \N__47426\,
            in2 => \_gnd_net_\,
            in3 => \N__47393\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47768\,
            in1 => \N__43232\,
            in2 => \_gnd_net_\,
            in3 => \N__47801\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44765\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__43236\,
            in1 => \N__47965\,
            in2 => \_gnd_net_\,
            in3 => \N__48005\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__44320\,
            in1 => \N__49409\,
            in2 => \_gnd_net_\,
            in3 => \N__44292\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49411\,
            in1 => \N__43406\,
            in2 => \_gnd_net_\,
            in3 => \N__43379\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43490\,
            in1 => \N__49412\,
            in2 => \_gnd_net_\,
            in3 => \N__43460\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49410\,
            in1 => \_gnd_net_\,
            in2 => \N__44390\,
            in3 => \N__44349\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43489\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49413\,
            in1 => \N__44461\,
            in2 => \N__50004\,
            in3 => \N__44421\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46861\,
            in1 => \N__43237\,
            in2 => \_gnd_net_\,
            in3 => \N__43619\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100111"
        )
    port map (
            in0 => \N__49106\,
            in1 => \N__45109\,
            in2 => \N__48787\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48157\,
            in1 => \N__44584\,
            in2 => \_gnd_net_\,
            in3 => \N__49104\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43093\,
            in3 => \N__43085\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52572\,
            ce => 'H',
            sr => \N__52231\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49105\,
            lcout => \current_shift_inst.N_1379_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__49107\,
            in1 => \N__45091\,
            in2 => \_gnd_net_\,
            in3 => \N__48760\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__45070\,
            in1 => \N__48730\,
            in2 => \_gnd_net_\,
            in3 => \N__49108\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48421\,
            in1 => \N__44779\,
            in2 => \_gnd_net_\,
            in3 => \N__49117\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50054\,
            in1 => \N__49501\,
            in2 => \N__43501\,
            in3 => \N__43468\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48658\,
            in1 => \N__45010\,
            in2 => \_gnd_net_\,
            in3 => \N__49119\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__49120\,
            in1 => \N__44986\,
            in2 => \_gnd_net_\,
            in3 => \N__48634\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49499\,
            in1 => \N__50055\,
            in2 => \N__46863\,
            in3 => \N__43620\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__49118\,
            in1 => \N__45055\,
            in2 => \_gnd_net_\,
            in3 => \N__48709\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48799\,
            in1 => \N__45130\,
            in2 => \_gnd_net_\,
            in3 => \N__49121\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50053\,
            in1 => \N__49500\,
            in2 => \N__43419\,
            in3 => \N__43380\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50061\,
            in1 => \N__49503\,
            in2 => \N__44770\,
            in3 => \N__44731\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__48919\,
            in1 => \N__45214\,
            in2 => \_gnd_net_\,
            in3 => \N__49165\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43500\,
            in1 => \N__49507\,
            in2 => \N__50100\,
            in3 => \N__43467\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49506\,
            in1 => \N__50056\,
            in2 => \N__44395\,
            in3 => \N__44353\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44324\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49504\,
            in1 => \N__50062\,
            in2 => \N__44329\,
            in3 => \N__44296\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__49166\,
            in1 => \N__48892\,
            in2 => \_gnd_net_\,
            in3 => \N__45196\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49505\,
            in1 => \N__50057\,
            in2 => \N__43420\,
            in3 => \N__43381\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43357\,
            in1 => \N__43345\,
            in2 => \N__43339\,
            in3 => \N__43324\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__43621\,
            in1 => \N__50066\,
            in2 => \N__46867\,
            in3 => \N__49502\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43848\,
            in1 => \N__43597\,
            in2 => \_gnd_net_\,
            in3 => \N__50536\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => \elapsed_time_ns_1_RNIJ53T9_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43591\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43578\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45330\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43543\,
            in1 => \N__46942\,
            in2 => \_gnd_net_\,
            in3 => \N__50538\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43537\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43525\,
            in1 => \N__43882\,
            in2 => \_gnd_net_\,
            in3 => \N__50537\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43519\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50532\,
            in1 => \N__43687\,
            in2 => \_gnd_net_\,
            in3 => \N__46180\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => \elapsed_time_ns_1_RNITUBN9_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43681\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__43657\,
            in1 => \_gnd_net_\,
            in2 => \N__50546\,
            in3 => \N__46264\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43821\,
            in1 => \N__43672\,
            in2 => \_gnd_net_\,
            in3 => \N__50530\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43666\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43656\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50531\,
            in1 => \N__43642\,
            in2 => \_gnd_net_\,
            in3 => \N__46228\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => \elapsed_time_ns_1_RNIL73T9_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43636\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43737\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43753\,
            in1 => \N__46279\,
            in2 => \_gnd_net_\,
            in3 => \N__50518\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50515\,
            in1 => \N__43783\,
            in2 => \_gnd_net_\,
            in3 => \N__43864\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43777\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50516\,
            in1 => \N__43768\,
            in2 => \_gnd_net_\,
            in3 => \N__46213\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43762\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43752\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43738\,
            in1 => \N__46198\,
            in2 => \_gnd_net_\,
            in3 => \N__50517\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45315\,
            in2 => \N__45651\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45624\,
            in2 => \N__45684\,
            in3 => \N__43690\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45603\,
            in2 => \N__45652\,
            in3 => \N__43867\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45625\,
            in2 => \N__45573\,
            in3 => \N__43852\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45543\,
            in2 => \N__45604\,
            in3 => \N__43828\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45519\,
            in2 => \N__45574\,
            in3 => \N__43801\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45544\,
            in2 => \N__45492\,
            in3 => \N__43798\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45942\,
            in2 => \N__45523\,
            in3 => \N__43795\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__52637\,
            ce => \N__43972\,
            sr => \N__52173\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45493\,
            in2 => \N__45909\,
            in3 => \N__43792\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45882\,
            in2 => \N__45946\,
            in3 => \N__43789\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45855\,
            in2 => \N__45910\,
            in3 => \N__43786\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45883\,
            in2 => \N__45829\,
            in3 => \N__43909\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45798\,
            in2 => \N__45859\,
            in3 => \N__43906\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45825\,
            in2 => \N__45777\,
            in3 => \N__43903\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45799\,
            in2 => \N__45747\,
            in3 => \N__43900\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45711\,
            in2 => \N__45778\,
            in3 => \N__43897\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__52631\,
            ce => \N__43970\,
            sr => \N__52175\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46164\,
            in2 => \N__45751\,
            in3 => \N__43894\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46140\,
            in2 => \N__45718\,
            in3 => \N__43891\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46165\,
            in2 => \N__46119\,
            in3 => \N__43888\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46141\,
            in2 => \N__46093\,
            in3 => \N__43885\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46062\,
            in2 => \N__46120\,
            in3 => \N__43999\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46089\,
            in2 => \N__46041\,
            in3 => \N__43996\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46063\,
            in2 => \N__46011\,
            in3 => \N__43993\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45972\,
            in2 => \N__46042\,
            in3 => \N__43990\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__52625\,
            ce => \N__43963\,
            sr => \N__52177\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46392\,
            in2 => \N__46015\,
            in3 => \N__43987\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__52619\,
            ce => \N__43971\,
            sr => \N__52182\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46362\,
            in2 => \N__45979\,
            in3 => \N__43984\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__52619\,
            ce => \N__43971\,
            sr => \N__52182\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46336\,
            in2 => \N__46396\,
            in3 => \N__43981\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__52619\,
            ce => \N__43971\,
            sr => \N__52182\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46312\,
            in2 => \N__46366\,
            in3 => \N__43978\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__52619\,
            ce => \N__43971\,
            sr => \N__52182\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43975\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52619\,
            ce => \N__43971\,
            sr => \N__52182\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49352\,
            in1 => \N__50082\,
            in2 => \N__44062\,
            in3 => \N__44022\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47858\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49351\,
            in1 => \N__50081\,
            in2 => \N__47299\,
            in3 => \N__47319\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50083\,
            in1 => \N__49353\,
            in2 => \N__47107\,
            in3 => \N__47127\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49349\,
            in1 => \N__50080\,
            in2 => \N__47644\,
            in3 => \N__47664\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__50078\,
            in1 => \N__49348\,
            in2 => \N__48360\,
            in3 => \N__48393\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__49350\,
            in1 => \N__47036\,
            in2 => \N__47074\,
            in3 => \N__50079\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__50084\,
            in1 => \N__49354\,
            in2 => \N__47401\,
            in3 => \N__47434\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49333\,
            in1 => \N__44272\,
            in2 => \N__50085\,
            in3 => \N__44247\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__44271\,
            in1 => \N__49332\,
            in2 => \N__44248\,
            in3 => \N__49997\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44226\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52600\,
            ce => \N__44195\,
            sr => \N__52193\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__44148\,
            in1 => \N__49998\,
            in2 => \N__44170\,
            in3 => \N__49331\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__49999\,
            in1 => \N__44166\,
            in2 => \N__49408\,
            in3 => \N__44147\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__44086\,
            in1 => \N__44095\,
            in2 => \_gnd_net_\,
            in3 => \N__49327\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44119\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49326\,
            in2 => \N__44089\,
            in3 => \N__44085\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49367\,
            in1 => \N__50012\,
            in2 => \N__48070\,
            in3 => \N__48032\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50006\,
            in1 => \N__49364\,
            in2 => \N__44061\,
            in3 => \N__44026\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__49368\,
            in1 => \N__50007\,
            in2 => \N__44548\,
            in3 => \N__44575\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__44574\,
            in1 => \N__44543\,
            in2 => \N__50086\,
            in3 => \N__49369\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49370\,
            in1 => \N__50013\,
            in2 => \N__48010\,
            in3 => \N__47960\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50014\,
            in1 => \N__49366\,
            in2 => \N__47910\,
            in3 => \N__47934\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49363\,
            in1 => \N__50005\,
            in2 => \N__44527\,
            in3 => \N__44484\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__50011\,
            in1 => \N__49365\,
            in2 => \N__47731\,
            in3 => \N__47694\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__44460\,
            in1 => \N__49465\,
            in2 => \N__44425\,
            in3 => \N__49824\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49471\,
            in1 => \N__44391\,
            in2 => \N__50000\,
            in3 => \N__44348\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__47806\,
            in1 => \N__49817\,
            in2 => \N__47775\,
            in3 => \N__49468\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49470\,
            in1 => \N__44328\,
            in2 => \N__50003\,
            in3 => \N__44291\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__44761\,
            in1 => \N__49469\,
            in2 => \N__44730\,
            in3 => \N__49825\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49467\,
            in1 => \N__44683\,
            in2 => \N__50001\,
            in3 => \N__44655\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \N__50755\,
            in1 => \N__49472\,
            in2 => \N__44705\,
            in3 => \N__49829\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49466\,
            in1 => \N__44682\,
            in2 => \N__50002\,
            in3 => \N__44656\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44635\,
            in2 => \N__50676\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48206\,
            in2 => \N__44626\,
            in3 => \N__50749\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__50750\,
            in1 => \N__49680\,
            in2 => \N__44608\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44593\,
            in2 => \N__49884\,
            in3 => \N__44578\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49684\,
            in2 => \N__44953\,
            in3 => \N__44932\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44929\,
            in2 => \N__49885\,
            in3 => \N__44905\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49688\,
            in2 => \N__46753\,
            in3 => \N__44890\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49689\,
            in2 => \N__48286\,
            in3 => \N__44875\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49706\,
            in2 => \N__44872\,
            in3 => \N__44845\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44842\,
            in2 => \N__49890\,
            in3 => \N__44821\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49710\,
            in2 => \N__44818\,
            in3 => \N__44791\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44788\,
            in2 => \N__49891\,
            in3 => \N__44773\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49714\,
            in2 => \N__45121\,
            in3 => \N__45103\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45100\,
            in2 => \N__49892\,
            in3 => \N__45085\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49718\,
            in2 => \N__45082\,
            in3 => \N__45064\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45061\,
            in2 => \N__49893\,
            in3 => \N__45049\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49894\,
            in2 => \N__45046\,
            in3 => \N__45025\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45022\,
            in2 => \N__50046\,
            in3 => \N__45004\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49898\,
            in2 => \N__45001\,
            in3 => \N__44980\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44977\,
            in2 => \N__50047\,
            in3 => \N__44956\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49902\,
            in2 => \N__45289\,
            in3 => \N__45262\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45259\,
            in2 => \N__50048\,
            in3 => \N__45235\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49906\,
            in2 => \N__45232\,
            in3 => \N__45208\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45205\,
            in2 => \N__50049\,
            in3 => \N__45190\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49910\,
            in2 => \N__45187\,
            in3 => \N__45169\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45166\,
            in2 => \N__50050\,
            in3 => \N__45151\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49914\,
            in2 => \N__45148\,
            in3 => \N__45139\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45136\,
            in2 => \N__50051\,
            in3 => \N__45124\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49918\,
            in2 => \N__45463\,
            in3 => \N__45439\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45436\,
            in2 => \N__50052\,
            in3 => \N__45421\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49922\,
            in2 => \N__45418\,
            in3 => \N__45388\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__45385\,
            in1 => \N__49195\,
            in2 => \N__49177\,
            in3 => \N__45370\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45355\,
            in1 => \N__46600\,
            in2 => \_gnd_net_\,
            in3 => \N__50540\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => \elapsed_time_ns_1_RNI58DN9_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45349\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50539\,
            in1 => \N__45331\,
            in2 => \_gnd_net_\,
            in3 => \N__46297\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46522\,
            in1 => \N__45303\,
            in2 => \_gnd_net_\,
            in3 => \N__45292\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46461\,
            in1 => \N__45677\,
            in2 => \_gnd_net_\,
            in3 => \N__45655\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46523\,
            in1 => \N__45644\,
            in2 => \_gnd_net_\,
            in3 => \N__45628\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46462\,
            in1 => \N__45623\,
            in2 => \_gnd_net_\,
            in3 => \N__45607\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46524\,
            in1 => \N__45596\,
            in2 => \_gnd_net_\,
            in3 => \N__45577\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46463\,
            in1 => \N__45561\,
            in2 => \_gnd_net_\,
            in3 => \N__45547\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46525\,
            in1 => \N__45542\,
            in2 => \_gnd_net_\,
            in3 => \N__45526\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46464\,
            in1 => \N__45512\,
            in2 => \_gnd_net_\,
            in3 => \N__45496\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__52657\,
            ce => \N__47469\,
            sr => \N__52169\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46460\,
            in1 => \N__45485\,
            in2 => \_gnd_net_\,
            in3 => \N__45466\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46508\,
            in1 => \N__45941\,
            in2 => \_gnd_net_\,
            in3 => \N__45913\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46457\,
            in1 => \N__45902\,
            in2 => \_gnd_net_\,
            in3 => \N__45886\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46505\,
            in1 => \N__45876\,
            in2 => \_gnd_net_\,
            in3 => \N__45862\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46458\,
            in1 => \N__45848\,
            in2 => \_gnd_net_\,
            in3 => \N__45832\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46506\,
            in1 => \N__45821\,
            in2 => \_gnd_net_\,
            in3 => \N__45802\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46459\,
            in1 => \N__45797\,
            in2 => \_gnd_net_\,
            in3 => \N__45781\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46507\,
            in1 => \N__45770\,
            in2 => \_gnd_net_\,
            in3 => \N__45754\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__52655\,
            ce => \N__47470\,
            sr => \N__52170\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46501\,
            in1 => \N__45740\,
            in2 => \_gnd_net_\,
            in3 => \N__45721\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46518\,
            in1 => \N__45710\,
            in2 => \_gnd_net_\,
            in3 => \N__45688\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46502\,
            in1 => \N__46158\,
            in2 => \_gnd_net_\,
            in3 => \N__46144\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46519\,
            in1 => \N__46139\,
            in2 => \_gnd_net_\,
            in3 => \N__46123\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46503\,
            in1 => \N__46112\,
            in2 => \_gnd_net_\,
            in3 => \N__46096\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46520\,
            in1 => \N__46085\,
            in2 => \_gnd_net_\,
            in3 => \N__46066\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46504\,
            in1 => \N__46061\,
            in2 => \_gnd_net_\,
            in3 => \N__46045\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46521\,
            in1 => \N__46034\,
            in2 => \_gnd_net_\,
            in3 => \N__46018\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__52649\,
            ce => \N__47468\,
            sr => \N__52171\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46465\,
            in1 => \N__46010\,
            in2 => \_gnd_net_\,
            in3 => \N__45982\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__52642\,
            ce => \N__47467\,
            sr => \N__52172\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46499\,
            in1 => \N__45971\,
            in2 => \_gnd_net_\,
            in3 => \N__45949\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__52642\,
            ce => \N__47467\,
            sr => \N__52172\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46466\,
            in1 => \N__46385\,
            in2 => \_gnd_net_\,
            in3 => \N__46369\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__52642\,
            ce => \N__47467\,
            sr => \N__52172\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46500\,
            in1 => \N__46355\,
            in2 => \_gnd_net_\,
            in3 => \N__46339\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__52642\,
            ce => \N__47467\,
            sr => \N__52172\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46467\,
            in1 => \N__46332\,
            in2 => \_gnd_net_\,
            in3 => \N__46318\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__52642\,
            ce => \N__47467\,
            sr => \N__52172\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__46311\,
            in1 => \N__46468\,
            in2 => \_gnd_net_\,
            in3 => \N__46315\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52642\,
            ce => \N__47467\,
            sr => \N__52172\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46612\,
            in1 => \N__50619\,
            in2 => \_gnd_net_\,
            in3 => \N__50524\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46290\,
            in1 => \N__46275\,
            in2 => \N__46263\,
            in3 => \N__46557\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46246\,
            in1 => \N__46627\,
            in2 => \_gnd_net_\,
            in3 => \N__50525\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46240\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46224\,
            in1 => \N__46209\,
            in2 => \N__46197\,
            in3 => \N__46176\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50559\,
            in2 => \N__46705\,
            in3 => \N__49023\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__46698\,
            in1 => \N__46873\,
            in2 => \N__46681\,
            in3 => \N__46678\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46647\,
            in2 => \N__46666\,
            in3 => \N__46663\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46623\,
            in1 => \N__46611\,
            in2 => \N__46599\,
            in3 => \N__46569\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46546\,
            in1 => \N__46558\,
            in2 => \_gnd_net_\,
            in3 => \N__50477\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46540\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46908\,
            in1 => \N__47605\,
            in2 => \_gnd_net_\,
            in3 => \N__50478\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47535\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46989\,
            in1 => \N__46971\,
            in2 => \N__50592\,
            in3 => \N__46953\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46938\,
            in1 => \N__46920\,
            in2 => \N__46909\,
            in3 => \N__46737\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46894\,
            in1 => \N__46888\,
            in2 => \N__46882\,
            in3 => \N__46879\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46862\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__46771\,
            in1 => \N__49415\,
            in2 => \N__46804\,
            in3 => \N__50096\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49414\,
            in1 => \N__46803\,
            in2 => \N__50105\,
            in3 => \N__46770\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46726\,
            in1 => \N__46738\,
            in2 => \_gnd_net_\,
            in3 => \N__50526\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46720\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47604\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__47581\,
            in1 => \N__47539\,
            in2 => \_gnd_net_\,
            in3 => \N__47506\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__47433\,
            in1 => \N__49380\,
            in2 => \N__47400\,
            in3 => \N__50075\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__50269\,
            in1 => \N__50244\,
            in2 => \_gnd_net_\,
            in3 => \N__50300\,
            lcout => \current_shift_inst.timer_s1.N_164_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__47320\,
            in1 => \N__50073\,
            in2 => \N__47298\,
            in3 => \N__49378\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50243\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__47131\,
            in1 => \N__50074\,
            in2 => \N__47106\,
            in3 => \N__49379\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49377\,
            in1 => \N__47070\,
            in2 => \N__50104\,
            in3 => \N__47038\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50248\,
            in2 => \_gnd_net_\,
            in3 => \N__50302\,
            lcout => \current_shift_inst.timer_s1.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49371\,
            in1 => \N__48121\,
            in2 => \N__50091\,
            in3 => \N__48096\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__48066\,
            in1 => \N__49375\,
            in2 => \N__48037\,
            in3 => \N__50032\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49376\,
            in1 => \N__48006\,
            in2 => \N__50092\,
            in3 => \N__47964\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__47938\,
            in1 => \N__50037\,
            in2 => \N__47914\,
            in3 => \N__49372\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49373\,
            in1 => \N__47867\,
            in2 => \N__50090\,
            in3 => \N__47829\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__47802\,
            in1 => \N__50033\,
            in2 => \N__47776\,
            in3 => \N__49374\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49347\,
            in1 => \N__47727\,
            in2 => \N__50089\,
            in3 => \N__47698\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__49360\,
            in1 => \N__50018\,
            in2 => \N__47671\,
            in3 => \N__47640\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__49346\,
            in1 => \N__48394\,
            in2 => \N__50087\,
            in3 => \N__48361\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__49345\,
            in1 => \N__48334\,
            in2 => \N__48313\,
            in3 => \N__48213\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__49361\,
            in1 => \N__50019\,
            in2 => \N__48253\,
            in3 => \N__48273\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__48274\,
            in1 => \N__48249\,
            in2 => \N__50088\,
            in3 => \N__49362\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50694\,
            in2 => \N__50677\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48205\,
            in2 => \N__48184\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48175\,
            in2 => \N__49881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49671\,
            in2 => \N__48166\,
            in3 => \N__48145\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48142\,
            in2 => \N__49882\,
            in3 => \N__48124\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49675\,
            in2 => \N__48589\,
            in3 => \N__48565\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48562\,
            in2 => \N__49883\,
            in3 => \N__48541\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49679\,
            in2 => \N__48538\,
            in3 => \N__48517\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49690\,
            in2 => \N__48514\,
            in3 => \N__48487\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48484\,
            in2 => \N__49886\,
            in3 => \N__48460\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49694\,
            in2 => \N__48457\,
            in3 => \N__48433\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48430\,
            in2 => \N__49887\,
            in3 => \N__48409\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49698\,
            in2 => \N__48406\,
            in3 => \N__48772\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48769\,
            in2 => \N__49888\,
            in3 => \N__48748\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49702\,
            in2 => \N__48745\,
            in3 => \N__48718\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48715\,
            in2 => \N__49889\,
            in3 => \N__48697\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48694\,
            in2 => \N__49947\,
            in3 => \N__48673\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49767\,
            in2 => \N__48670\,
            in3 => \N__48646\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48643\,
            in2 => \N__49948\,
            in3 => \N__48622\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49771\,
            in2 => \N__48619\,
            in3 => \N__48592\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48982\,
            in2 => \N__49949\,
            in3 => \N__48958\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49775\,
            in2 => \N__48955\,
            in3 => \N__48931\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48928\,
            in2 => \N__49950\,
            in3 => \N__48907\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49779\,
            in2 => \N__48904\,
            in3 => \N__48880\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49951\,
            in2 => \N__48877\,
            in3 => \N__48853\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48850\,
            in2 => \N__50067\,
            in3 => \N__48829\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49955\,
            in2 => \N__48826\,
            in3 => \N__48814\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48811\,
            in2 => \N__50068\,
            in3 => \N__48790\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49959\,
            in2 => \N__50191\,
            in3 => \N__50167\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50164\,
            in2 => \N__50069\,
            in3 => \N__50143\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49963\,
            in2 => \N__50140\,
            in3 => \N__50116\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__49964\,
            in1 => \N__49495\,
            in2 => \_gnd_net_\,
            in3 => \N__49198\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__49189\,
            in1 => \N__49183\,
            in2 => \_gnd_net_\,
            in3 => \N__49173\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49030\,
            in1 => \N__49012\,
            in2 => \_gnd_net_\,
            in3 => \N__50527\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49006\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50379\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50574\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__50620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50575\,
            in1 => \N__50596\,
            in2 => \_gnd_net_\,
            in3 => \N__50523\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50380\,
            in1 => \N__50563\,
            in2 => \_gnd_net_\,
            in3 => \N__50522\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50342\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52632\,
            ce => 'H',
            sr => \N__52183\
        );

    \current_shift_inst.start_timer_s1_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__50357\,
            in1 => \N__50266\,
            in2 => \_gnd_net_\,
            in3 => \N__50344\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52632\,
            ce => 'H',
            sr => \N__52183\
        );

    \current_shift_inst.stop_timer_s1_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__50358\,
            in1 => \N__50343\,
            in2 => \N__50301\,
            in3 => \N__50267\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52632\,
            ce => 'H',
            sr => \N__52183\
        );

    \current_shift_inst.timer_s1.running_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__50296\,
            in1 => \N__50239\,
            in2 => \_gnd_net_\,
            in3 => \N__50268\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52632\,
            ce => 'H',
            sr => \N__52183\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50217\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52620\,
            ce => 'H',
            sr => \N__52194\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51667\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52620\,
            ce => 'H',
            sr => \N__52194\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__51475\,
            in1 => \N__50748\,
            in2 => \_gnd_net_\,
            in3 => \N__50698\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53051\,
            in2 => \_gnd_net_\,
            in3 => \N__51704\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__52757\,
            in1 => \N__51903\,
            in2 => \N__50650\,
            in3 => \N__53175\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__50646\,
            in1 => \N__52700\,
            in2 => \_gnd_net_\,
            in3 => \N__52874\,
            lcout => \current_shift_inst.PI_CTRL.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53052\,
            in1 => \N__50635\,
            in2 => \N__51711\,
            in3 => \N__52770\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__50647\,
            in1 => \N__52876\,
            in2 => \N__52718\,
            in3 => \N__53111\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__52875\,
            in1 => \N__50645\,
            in2 => \N__53113\,
            in3 => \N__52701\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51890\,
            in2 => \_gnd_net_\,
            in3 => \N__53168\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__52900\,
            in1 => \N__53124\,
            in2 => \N__51958\,
            in3 => \N__52823\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__52983\,
            in1 => \N__51967\,
            in2 => \N__51961\,
            in3 => \N__52938\,
            lcout => \current_shift_inst.PI_CTRL.N_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53104\,
            in2 => \_gnd_net_\,
            in3 => \N__52976\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_i_LC_24_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__51945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__52834\,
            in1 => \N__52918\,
            in2 => \N__52728\,
            in3 => \N__51904\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52650\,
            ce => 'H',
            sr => \N__52217\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52916\,
            lcout => pwm_duty_input_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52650\,
            ce => 'H',
            sr => \N__52217\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51769\,
            in2 => \_gnd_net_\,
            in3 => \N__53004\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52650\,
            ce => 'H',
            sr => \N__52217\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51742\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52650\,
            ce => 'H',
            sr => \N__52217\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__52917\,
            in1 => \N__52833\,
            in2 => \N__51715\,
            in3 => \N__52722\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52650\,
            ce => 'H',
            sr => \N__52217\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__52920\,
            in1 => \N__52830\,
            in2 => \N__53182\,
            in3 => \N__52726\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52643\,
            ce => 'H',
            sr => \N__52223\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__52832\,
            in1 => \N__53140\,
            in2 => \N__53131\,
            in3 => \N__53112\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52643\,
            ce => 'H',
            sr => \N__52223\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__52831\,
            in1 => \N__52921\,
            in2 => \N__52729\,
            in3 => \N__53056\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52643\,
            ce => 'H',
            sr => \N__52223\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53003\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52643\,
            ce => 'H',
            sr => \N__52223\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__52984\,
            in1 => \N__52948\,
            in2 => \_gnd_net_\,
            in3 => \N__52942\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52643\,
            ce => 'H',
            sr => \N__52223\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__52919\,
            in1 => \N__52829\,
            in2 => \N__52774\,
            in3 => \N__52727\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52638\,
            ce => 'H',
            sr => \N__52232\
        );
end \INTERFACE\;
