// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 23 2024 20:10:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    error_pin,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    input error_pin;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__53076;
    wire N__53075;
    wire N__53074;
    wire N__53065;
    wire N__53064;
    wire N__53063;
    wire N__53056;
    wire N__53055;
    wire N__53054;
    wire N__53047;
    wire N__53046;
    wire N__53045;
    wire N__53038;
    wire N__53037;
    wire N__53036;
    wire N__53029;
    wire N__53028;
    wire N__53027;
    wire N__53020;
    wire N__53019;
    wire N__53018;
    wire N__53011;
    wire N__53010;
    wire N__53009;
    wire N__53002;
    wire N__53001;
    wire N__53000;
    wire N__52993;
    wire N__52992;
    wire N__52991;
    wire N__52984;
    wire N__52983;
    wire N__52982;
    wire N__52975;
    wire N__52974;
    wire N__52973;
    wire N__52966;
    wire N__52965;
    wire N__52964;
    wire N__52947;
    wire N__52944;
    wire N__52941;
    wire N__52940;
    wire N__52939;
    wire N__52936;
    wire N__52933;
    wire N__52930;
    wire N__52929;
    wire N__52926;
    wire N__52921;
    wire N__52918;
    wire N__52915;
    wire N__52910;
    wire N__52905;
    wire N__52902;
    wire N__52899;
    wire N__52896;
    wire N__52895;
    wire N__52892;
    wire N__52889;
    wire N__52886;
    wire N__52883;
    wire N__52878;
    wire N__52875;
    wire N__52872;
    wire N__52869;
    wire N__52866;
    wire N__52863;
    wire N__52862;
    wire N__52861;
    wire N__52858;
    wire N__52853;
    wire N__52848;
    wire N__52845;
    wire N__52842;
    wire N__52839;
    wire N__52836;
    wire N__52833;
    wire N__52830;
    wire N__52827;
    wire N__52826;
    wire N__52825;
    wire N__52822;
    wire N__52819;
    wire N__52816;
    wire N__52813;
    wire N__52810;
    wire N__52807;
    wire N__52804;
    wire N__52799;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52781;
    wire N__52778;
    wire N__52775;
    wire N__52774;
    wire N__52771;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52757;
    wire N__52754;
    wire N__52751;
    wire N__52746;
    wire N__52743;
    wire N__52740;
    wire N__52737;
    wire N__52734;
    wire N__52731;
    wire N__52728;
    wire N__52727;
    wire N__52726;
    wire N__52723;
    wire N__52720;
    wire N__52717;
    wire N__52710;
    wire N__52707;
    wire N__52704;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52692;
    wire N__52691;
    wire N__52690;
    wire N__52689;
    wire N__52688;
    wire N__52687;
    wire N__52684;
    wire N__52673;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52649;
    wire N__52648;
    wire N__52647;
    wire N__52646;
    wire N__52635;
    wire N__52634;
    wire N__52631;
    wire N__52628;
    wire N__52627;
    wire N__52626;
    wire N__52625;
    wire N__52624;
    wire N__52621;
    wire N__52618;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52593;
    wire N__52590;
    wire N__52589;
    wire N__52588;
    wire N__52587;
    wire N__52586;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52566;
    wire N__52563;
    wire N__52562;
    wire N__52561;
    wire N__52560;
    wire N__52557;
    wire N__52552;
    wire N__52549;
    wire N__52542;
    wire N__52539;
    wire N__52536;
    wire N__52533;
    wire N__52532;
    wire N__52531;
    wire N__52528;
    wire N__52523;
    wire N__52518;
    wire N__52515;
    wire N__52512;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52500;
    wire N__52499;
    wire N__52498;
    wire N__52497;
    wire N__52496;
    wire N__52495;
    wire N__52494;
    wire N__52493;
    wire N__52492;
    wire N__52491;
    wire N__52490;
    wire N__52489;
    wire N__52488;
    wire N__52487;
    wire N__52486;
    wire N__52485;
    wire N__52484;
    wire N__52483;
    wire N__52482;
    wire N__52481;
    wire N__52480;
    wire N__52479;
    wire N__52478;
    wire N__52477;
    wire N__52476;
    wire N__52475;
    wire N__52474;
    wire N__52473;
    wire N__52472;
    wire N__52471;
    wire N__52470;
    wire N__52469;
    wire N__52468;
    wire N__52467;
    wire N__52466;
    wire N__52465;
    wire N__52464;
    wire N__52463;
    wire N__52462;
    wire N__52461;
    wire N__52460;
    wire N__52459;
    wire N__52458;
    wire N__52457;
    wire N__52456;
    wire N__52455;
    wire N__52454;
    wire N__52453;
    wire N__52452;
    wire N__52451;
    wire N__52450;
    wire N__52449;
    wire N__52448;
    wire N__52447;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52443;
    wire N__52442;
    wire N__52441;
    wire N__52440;
    wire N__52439;
    wire N__52438;
    wire N__52437;
    wire N__52436;
    wire N__52435;
    wire N__52434;
    wire N__52433;
    wire N__52432;
    wire N__52431;
    wire N__52430;
    wire N__52429;
    wire N__52428;
    wire N__52427;
    wire N__52426;
    wire N__52425;
    wire N__52424;
    wire N__52423;
    wire N__52422;
    wire N__52421;
    wire N__52420;
    wire N__52419;
    wire N__52418;
    wire N__52417;
    wire N__52416;
    wire N__52415;
    wire N__52414;
    wire N__52413;
    wire N__52412;
    wire N__52411;
    wire N__52410;
    wire N__52409;
    wire N__52408;
    wire N__52407;
    wire N__52406;
    wire N__52405;
    wire N__52404;
    wire N__52403;
    wire N__52402;
    wire N__52401;
    wire N__52400;
    wire N__52399;
    wire N__52398;
    wire N__52397;
    wire N__52396;
    wire N__52395;
    wire N__52394;
    wire N__52393;
    wire N__52392;
    wire N__52391;
    wire N__52390;
    wire N__52389;
    wire N__52388;
    wire N__52387;
    wire N__52386;
    wire N__52385;
    wire N__52384;
    wire N__52383;
    wire N__52382;
    wire N__52381;
    wire N__52380;
    wire N__52379;
    wire N__52378;
    wire N__52377;
    wire N__52376;
    wire N__52375;
    wire N__52374;
    wire N__52373;
    wire N__52372;
    wire N__52371;
    wire N__52370;
    wire N__52369;
    wire N__52368;
    wire N__52367;
    wire N__52366;
    wire N__52365;
    wire N__52092;
    wire N__52089;
    wire N__52088;
    wire N__52087;
    wire N__52086;
    wire N__52085;
    wire N__52084;
    wire N__52083;
    wire N__52082;
    wire N__52079;
    wire N__52076;
    wire N__52073;
    wire N__52070;
    wire N__52067;
    wire N__52064;
    wire N__52061;
    wire N__52058;
    wire N__52055;
    wire N__52052;
    wire N__52049;
    wire N__52048;
    wire N__52047;
    wire N__52046;
    wire N__52045;
    wire N__52044;
    wire N__52043;
    wire N__52042;
    wire N__52041;
    wire N__52040;
    wire N__52039;
    wire N__52038;
    wire N__52037;
    wire N__52036;
    wire N__52035;
    wire N__52034;
    wire N__52033;
    wire N__52032;
    wire N__52031;
    wire N__52030;
    wire N__52027;
    wire N__52026;
    wire N__52025;
    wire N__52024;
    wire N__52023;
    wire N__52022;
    wire N__52021;
    wire N__52020;
    wire N__52019;
    wire N__52018;
    wire N__52017;
    wire N__52016;
    wire N__52015;
    wire N__52014;
    wire N__52013;
    wire N__52012;
    wire N__52011;
    wire N__52010;
    wire N__52009;
    wire N__52008;
    wire N__52007;
    wire N__52006;
    wire N__52005;
    wire N__52004;
    wire N__52003;
    wire N__52002;
    wire N__52001;
    wire N__52000;
    wire N__51999;
    wire N__51998;
    wire N__51997;
    wire N__51996;
    wire N__51995;
    wire N__51994;
    wire N__51993;
    wire N__51992;
    wire N__51991;
    wire N__51990;
    wire N__51989;
    wire N__51988;
    wire N__51987;
    wire N__51986;
    wire N__51983;
    wire N__51982;
    wire N__51981;
    wire N__51980;
    wire N__51979;
    wire N__51978;
    wire N__51977;
    wire N__51976;
    wire N__51975;
    wire N__51974;
    wire N__51973;
    wire N__51972;
    wire N__51971;
    wire N__51970;
    wire N__51969;
    wire N__51968;
    wire N__51967;
    wire N__51966;
    wire N__51965;
    wire N__51964;
    wire N__51963;
    wire N__51962;
    wire N__51961;
    wire N__51960;
    wire N__51959;
    wire N__51958;
    wire N__51957;
    wire N__51956;
    wire N__51955;
    wire N__51954;
    wire N__51953;
    wire N__51952;
    wire N__51951;
    wire N__51948;
    wire N__51947;
    wire N__51946;
    wire N__51945;
    wire N__51944;
    wire N__51943;
    wire N__51942;
    wire N__51941;
    wire N__51940;
    wire N__51939;
    wire N__51936;
    wire N__51935;
    wire N__51934;
    wire N__51933;
    wire N__51932;
    wire N__51929;
    wire N__51928;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51687;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51677;
    wire N__51676;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51660;
    wire N__51657;
    wire N__51654;
    wire N__51651;
    wire N__51648;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51627;
    wire N__51624;
    wire N__51621;
    wire N__51618;
    wire N__51615;
    wire N__51612;
    wire N__51609;
    wire N__51606;
    wire N__51605;
    wire N__51604;
    wire N__51597;
    wire N__51594;
    wire N__51591;
    wire N__51588;
    wire N__51585;
    wire N__51582;
    wire N__51579;
    wire N__51576;
    wire N__51573;
    wire N__51570;
    wire N__51567;
    wire N__51564;
    wire N__51563;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51545;
    wire N__51542;
    wire N__51539;
    wire N__51536;
    wire N__51533;
    wire N__51528;
    wire N__51527;
    wire N__51524;
    wire N__51521;
    wire N__51516;
    wire N__51513;
    wire N__51510;
    wire N__51507;
    wire N__51504;
    wire N__51501;
    wire N__51498;
    wire N__51497;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51474;
    wire N__51471;
    wire N__51468;
    wire N__51465;
    wire N__51462;
    wire N__51459;
    wire N__51456;
    wire N__51453;
    wire N__51450;
    wire N__51449;
    wire N__51446;
    wire N__51443;
    wire N__51440;
    wire N__51437;
    wire N__51434;
    wire N__51431;
    wire N__51426;
    wire N__51425;
    wire N__51422;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51405;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51393;
    wire N__51390;
    wire N__51387;
    wire N__51384;
    wire N__51381;
    wire N__51380;
    wire N__51379;
    wire N__51378;
    wire N__51375;
    wire N__51374;
    wire N__51371;
    wire N__51370;
    wire N__51369;
    wire N__51368;
    wire N__51367;
    wire N__51364;
    wire N__51361;
    wire N__51360;
    wire N__51359;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51346;
    wire N__51337;
    wire N__51328;
    wire N__51323;
    wire N__51320;
    wire N__51317;
    wire N__51314;
    wire N__51309;
    wire N__51300;
    wire N__51299;
    wire N__51296;
    wire N__51293;
    wire N__51290;
    wire N__51287;
    wire N__51284;
    wire N__51279;
    wire N__51276;
    wire N__51273;
    wire N__51270;
    wire N__51267;
    wire N__51264;
    wire N__51261;
    wire N__51260;
    wire N__51257;
    wire N__51254;
    wire N__51253;
    wire N__51250;
    wire N__51247;
    wire N__51244;
    wire N__51239;
    wire N__51234;
    wire N__51231;
    wire N__51228;
    wire N__51225;
    wire N__51222;
    wire N__51221;
    wire N__51218;
    wire N__51215;
    wire N__51212;
    wire N__51207;
    wire N__51204;
    wire N__51201;
    wire N__51198;
    wire N__51195;
    wire N__51192;
    wire N__51191;
    wire N__51190;
    wire N__51187;
    wire N__51184;
    wire N__51181;
    wire N__51178;
    wire N__51171;
    wire N__51168;
    wire N__51165;
    wire N__51162;
    wire N__51159;
    wire N__51156;
    wire N__51153;
    wire N__51150;
    wire N__51149;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51120;
    wire N__51117;
    wire N__51116;
    wire N__51115;
    wire N__51112;
    wire N__51109;
    wire N__51106;
    wire N__51103;
    wire N__51100;
    wire N__51093;
    wire N__51090;
    wire N__51087;
    wire N__51084;
    wire N__51081;
    wire N__51080;
    wire N__51077;
    wire N__51074;
    wire N__51071;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51042;
    wire N__51039;
    wire N__51036;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51018;
    wire N__51015;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51003;
    wire N__51000;
    wire N__50997;
    wire N__50994;
    wire N__50991;
    wire N__50988;
    wire N__50985;
    wire N__50982;
    wire N__50979;
    wire N__50976;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50964;
    wire N__50961;
    wire N__50958;
    wire N__50955;
    wire N__50952;
    wire N__50949;
    wire N__50946;
    wire N__50943;
    wire N__50940;
    wire N__50937;
    wire N__50934;
    wire N__50931;
    wire N__50928;
    wire N__50925;
    wire N__50922;
    wire N__50919;
    wire N__50916;
    wire N__50913;
    wire N__50910;
    wire N__50907;
    wire N__50904;
    wire N__50901;
    wire N__50898;
    wire N__50895;
    wire N__50892;
    wire N__50891;
    wire N__50888;
    wire N__50885;
    wire N__50880;
    wire N__50879;
    wire N__50878;
    wire N__50877;
    wire N__50876;
    wire N__50875;
    wire N__50874;
    wire N__50873;
    wire N__50870;
    wire N__50869;
    wire N__50866;
    wire N__50861;
    wire N__50856;
    wire N__50853;
    wire N__50852;
    wire N__50851;
    wire N__50850;
    wire N__50849;
    wire N__50848;
    wire N__50847;
    wire N__50846;
    wire N__50845;
    wire N__50838;
    wire N__50837;
    wire N__50836;
    wire N__50835;
    wire N__50834;
    wire N__50833;
    wire N__50826;
    wire N__50825;
    wire N__50824;
    wire N__50823;
    wire N__50822;
    wire N__50819;
    wire N__50818;
    wire N__50817;
    wire N__50816;
    wire N__50815;
    wire N__50804;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50788;
    wire N__50785;
    wire N__50780;
    wire N__50777;
    wire N__50768;
    wire N__50765;
    wire N__50756;
    wire N__50751;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50718;
    wire N__50715;
    wire N__50712;
    wire N__50709;
    wire N__50708;
    wire N__50705;
    wire N__50702;
    wire N__50697;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50684;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50662;
    wire N__50657;
    wire N__50654;
    wire N__50651;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50639;
    wire N__50636;
    wire N__50633;
    wire N__50628;
    wire N__50627;
    wire N__50624;
    wire N__50621;
    wire N__50618;
    wire N__50617;
    wire N__50612;
    wire N__50609;
    wire N__50606;
    wire N__50601;
    wire N__50598;
    wire N__50595;
    wire N__50594;
    wire N__50591;
    wire N__50588;
    wire N__50583;
    wire N__50582;
    wire N__50579;
    wire N__50576;
    wire N__50575;
    wire N__50574;
    wire N__50573;
    wire N__50570;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50558;
    wire N__50549;
    wire N__50546;
    wire N__50541;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50529;
    wire N__50526;
    wire N__50523;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50511;
    wire N__50508;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50484;
    wire N__50481;
    wire N__50478;
    wire N__50477;
    wire N__50474;
    wire N__50471;
    wire N__50466;
    wire N__50463;
    wire N__50460;
    wire N__50457;
    wire N__50454;
    wire N__50451;
    wire N__50448;
    wire N__50447;
    wire N__50444;
    wire N__50441;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50426;
    wire N__50423;
    wire N__50420;
    wire N__50415;
    wire N__50414;
    wire N__50411;
    wire N__50408;
    wire N__50403;
    wire N__50400;
    wire N__50397;
    wire N__50396;
    wire N__50393;
    wire N__50390;
    wire N__50385;
    wire N__50382;
    wire N__50379;
    wire N__50376;
    wire N__50373;
    wire N__50370;
    wire N__50369;
    wire N__50366;
    wire N__50363;
    wire N__50358;
    wire N__50355;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50343;
    wire N__50340;
    wire N__50337;
    wire N__50336;
    wire N__50333;
    wire N__50330;
    wire N__50325;
    wire N__50322;
    wire N__50321;
    wire N__50318;
    wire N__50315;
    wire N__50310;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50300;
    wire N__50297;
    wire N__50294;
    wire N__50289;
    wire N__50288;
    wire N__50285;
    wire N__50282;
    wire N__50277;
    wire N__50276;
    wire N__50273;
    wire N__50270;
    wire N__50267;
    wire N__50262;
    wire N__50259;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50247;
    wire N__50246;
    wire N__50243;
    wire N__50240;
    wire N__50235;
    wire N__50234;
    wire N__50229;
    wire N__50226;
    wire N__50225;
    wire N__50222;
    wire N__50219;
    wire N__50214;
    wire N__50213;
    wire N__50208;
    wire N__50205;
    wire N__50204;
    wire N__50201;
    wire N__50198;
    wire N__50193;
    wire N__50192;
    wire N__50187;
    wire N__50184;
    wire N__50183;
    wire N__50180;
    wire N__50177;
    wire N__50172;
    wire N__50171;
    wire N__50168;
    wire N__50165;
    wire N__50160;
    wire N__50157;
    wire N__50156;
    wire N__50155;
    wire N__50152;
    wire N__50149;
    wire N__50148;
    wire N__50147;
    wire N__50146;
    wire N__50145;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50135;
    wire N__50132;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50108;
    wire N__50105;
    wire N__50098;
    wire N__50095;
    wire N__50088;
    wire N__50085;
    wire N__50082;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50061;
    wire N__50058;
    wire N__50057;
    wire N__50054;
    wire N__50051;
    wire N__50048;
    wire N__50045;
    wire N__50040;
    wire N__50037;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50015;
    wire N__50012;
    wire N__50009;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49995;
    wire N__49992;
    wire N__49991;
    wire N__49986;
    wire N__49983;
    wire N__49982;
    wire N__49981;
    wire N__49976;
    wire N__49973;
    wire N__49970;
    wire N__49965;
    wire N__49964;
    wire N__49961;
    wire N__49958;
    wire N__49957;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49941;
    wire N__49938;
    wire N__49935;
    wire N__49932;
    wire N__49929;
    wire N__49926;
    wire N__49923;
    wire N__49920;
    wire N__49917;
    wire N__49916;
    wire N__49913;
    wire N__49910;
    wire N__49905;
    wire N__49904;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49890;
    wire N__49887;
    wire N__49884;
    wire N__49881;
    wire N__49880;
    wire N__49875;
    wire N__49872;
    wire N__49871;
    wire N__49866;
    wire N__49865;
    wire N__49862;
    wire N__49859;
    wire N__49856;
    wire N__49851;
    wire N__49850;
    wire N__49847;
    wire N__49844;
    wire N__49843;
    wire N__49838;
    wire N__49835;
    wire N__49832;
    wire N__49827;
    wire N__49826;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49790;
    wire N__49789;
    wire N__49784;
    wire N__49781;
    wire N__49778;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49766;
    wire N__49763;
    wire N__49760;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49734;
    wire N__49731;
    wire N__49728;
    wire N__49725;
    wire N__49722;
    wire N__49719;
    wire N__49716;
    wire N__49713;
    wire N__49710;
    wire N__49707;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49686;
    wire N__49683;
    wire N__49680;
    wire N__49677;
    wire N__49674;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49664;
    wire N__49661;
    wire N__49658;
    wire N__49653;
    wire N__49650;
    wire N__49647;
    wire N__49644;
    wire N__49641;
    wire N__49640;
    wire N__49637;
    wire N__49634;
    wire N__49631;
    wire N__49628;
    wire N__49623;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49611;
    wire N__49610;
    wire N__49607;
    wire N__49604;
    wire N__49599;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49589;
    wire N__49586;
    wire N__49583;
    wire N__49578;
    wire N__49577;
    wire N__49574;
    wire N__49571;
    wire N__49568;
    wire N__49565;
    wire N__49562;
    wire N__49557;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49536;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49509;
    wire N__49506;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49479;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49458;
    wire N__49455;
    wire N__49452;
    wire N__49449;
    wire N__49446;
    wire N__49443;
    wire N__49440;
    wire N__49437;
    wire N__49434;
    wire N__49431;
    wire N__49428;
    wire N__49425;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49404;
    wire N__49401;
    wire N__49398;
    wire N__49395;
    wire N__49392;
    wire N__49389;
    wire N__49386;
    wire N__49383;
    wire N__49382;
    wire N__49379;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49362;
    wire N__49359;
    wire N__49356;
    wire N__49355;
    wire N__49352;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49342;
    wire N__49335;
    wire N__49332;
    wire N__49329;
    wire N__49328;
    wire N__49325;
    wire N__49324;
    wire N__49321;
    wire N__49318;
    wire N__49315;
    wire N__49308;
    wire N__49305;
    wire N__49302;
    wire N__49301;
    wire N__49298;
    wire N__49297;
    wire N__49294;
    wire N__49291;
    wire N__49288;
    wire N__49281;
    wire N__49278;
    wire N__49275;
    wire N__49272;
    wire N__49271;
    wire N__49270;
    wire N__49267;
    wire N__49264;
    wire N__49261;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49247;
    wire N__49244;
    wire N__49243;
    wire N__49240;
    wire N__49237;
    wire N__49234;
    wire N__49227;
    wire N__49224;
    wire N__49221;
    wire N__49220;
    wire N__49219;
    wire N__49216;
    wire N__49213;
    wire N__49210;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49196;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49166;
    wire N__49165;
    wire N__49162;
    wire N__49159;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49107;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49097;
    wire N__49094;
    wire N__49091;
    wire N__49086;
    wire N__49083;
    wire N__49082;
    wire N__49081;
    wire N__49076;
    wire N__49073;
    wire N__49070;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49058;
    wire N__49055;
    wire N__49052;
    wire N__49049;
    wire N__49044;
    wire N__49041;
    wire N__49040;
    wire N__49039;
    wire N__49038;
    wire N__49037;
    wire N__49036;
    wire N__49035;
    wire N__49034;
    wire N__49033;
    wire N__49032;
    wire N__49031;
    wire N__49030;
    wire N__49029;
    wire N__49028;
    wire N__49027;
    wire N__49026;
    wire N__49025;
    wire N__49024;
    wire N__49023;
    wire N__49022;
    wire N__49021;
    wire N__49020;
    wire N__49019;
    wire N__49018;
    wire N__49017;
    wire N__49016;
    wire N__49015;
    wire N__49014;
    wire N__49013;
    wire N__49012;
    wire N__49003;
    wire N__48994;
    wire N__48985;
    wire N__48976;
    wire N__48971;
    wire N__48962;
    wire N__48953;
    wire N__48944;
    wire N__48937;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48917;
    wire N__48914;
    wire N__48911;
    wire N__48908;
    wire N__48903;
    wire N__48902;
    wire N__48899;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48889;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48876;
    wire N__48873;
    wire N__48870;
    wire N__48867;
    wire N__48864;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48850;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48834;
    wire N__48831;
    wire N__48828;
    wire N__48827;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48807;
    wire N__48804;
    wire N__48801;
    wire N__48798;
    wire N__48797;
    wire N__48794;
    wire N__48791;
    wire N__48788;
    wire N__48785;
    wire N__48784;
    wire N__48779;
    wire N__48776;
    wire N__48773;
    wire N__48768;
    wire N__48765;
    wire N__48764;
    wire N__48761;
    wire N__48758;
    wire N__48755;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48740;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48728;
    wire N__48725;
    wire N__48722;
    wire N__48721;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48705;
    wire N__48702;
    wire N__48701;
    wire N__48698;
    wire N__48695;
    wire N__48694;
    wire N__48689;
    wire N__48686;
    wire N__48683;
    wire N__48678;
    wire N__48675;
    wire N__48674;
    wire N__48673;
    wire N__48668;
    wire N__48665;
    wire N__48662;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48650;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48635;
    wire N__48630;
    wire N__48627;
    wire N__48626;
    wire N__48623;
    wire N__48620;
    wire N__48619;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48603;
    wire N__48600;
    wire N__48599;
    wire N__48598;
    wire N__48593;
    wire N__48590;
    wire N__48587;
    wire N__48582;
    wire N__48579;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48567;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48557;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48543;
    wire N__48542;
    wire N__48541;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48519;
    wire N__48516;
    wire N__48513;
    wire N__48512;
    wire N__48509;
    wire N__48506;
    wire N__48505;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48489;
    wire N__48486;
    wire N__48485;
    wire N__48480;
    wire N__48479;
    wire N__48476;
    wire N__48473;
    wire N__48470;
    wire N__48465;
    wire N__48462;
    wire N__48461;
    wire N__48456;
    wire N__48455;
    wire N__48452;
    wire N__48449;
    wire N__48446;
    wire N__48441;
    wire N__48438;
    wire N__48437;
    wire N__48434;
    wire N__48431;
    wire N__48426;
    wire N__48425;
    wire N__48422;
    wire N__48419;
    wire N__48416;
    wire N__48411;
    wire N__48408;
    wire N__48407;
    wire N__48404;
    wire N__48401;
    wire N__48396;
    wire N__48395;
    wire N__48392;
    wire N__48389;
    wire N__48386;
    wire N__48381;
    wire N__48378;
    wire N__48377;
    wire N__48372;
    wire N__48371;
    wire N__48368;
    wire N__48365;
    wire N__48362;
    wire N__48357;
    wire N__48354;
    wire N__48353;
    wire N__48348;
    wire N__48347;
    wire N__48344;
    wire N__48341;
    wire N__48338;
    wire N__48333;
    wire N__48330;
    wire N__48327;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48314;
    wire N__48309;
    wire N__48306;
    wire N__48303;
    wire N__48300;
    wire N__48299;
    wire N__48298;
    wire N__48293;
    wire N__48290;
    wire N__48287;
    wire N__48282;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48261;
    wire N__48258;
    wire N__48257;
    wire N__48254;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48239;
    wire N__48234;
    wire N__48231;
    wire N__48230;
    wire N__48227;
    wire N__48224;
    wire N__48221;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48211;
    wire N__48206;
    wire N__48201;
    wire N__48198;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48186;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48171;
    wire N__48168;
    wire N__48167;
    wire N__48164;
    wire N__48161;
    wire N__48158;
    wire N__48155;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48126;
    wire N__48123;
    wire N__48122;
    wire N__48119;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48105;
    wire N__48104;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48080;
    wire N__48077;
    wire N__48074;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48047;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47975;
    wire N__47972;
    wire N__47969;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47910;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47871;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47861;
    wire N__47858;
    wire N__47855;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47840;
    wire N__47837;
    wire N__47834;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47822;
    wire N__47819;
    wire N__47816;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47726;
    wire N__47723;
    wire N__47720;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47688;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47676;
    wire N__47673;
    wire N__47670;
    wire N__47667;
    wire N__47664;
    wire N__47661;
    wire N__47660;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47643;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47600;
    wire N__47595;
    wire N__47586;
    wire N__47583;
    wire N__47580;
    wire N__47577;
    wire N__47574;
    wire N__47573;
    wire N__47570;
    wire N__47567;
    wire N__47562;
    wire N__47559;
    wire N__47556;
    wire N__47553;
    wire N__47550;
    wire N__47547;
    wire N__47544;
    wire N__47541;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47529;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47510;
    wire N__47507;
    wire N__47504;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47435;
    wire N__47432;
    wire N__47429;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47412;
    wire N__47411;
    wire N__47408;
    wire N__47405;
    wire N__47400;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47364;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47282;
    wire N__47279;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47210;
    wire N__47207;
    wire N__47204;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47181;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47153;
    wire N__47150;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47120;
    wire N__47115;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47091;
    wire N__47088;
    wire N__47085;
    wire N__47082;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47070;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47057;
    wire N__47054;
    wire N__47051;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47033;
    wire N__47030;
    wire N__47027;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46989;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46967;
    wire N__46964;
    wire N__46961;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46941;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46890;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46875;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46849;
    wire N__46848;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46842;
    wire N__46841;
    wire N__46840;
    wire N__46839;
    wire N__46838;
    wire N__46837;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46829;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46799;
    wire N__46790;
    wire N__46787;
    wire N__46784;
    wire N__46781;
    wire N__46778;
    wire N__46775;
    wire N__46772;
    wire N__46771;
    wire N__46770;
    wire N__46769;
    wire N__46768;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46764;
    wire N__46763;
    wire N__46762;
    wire N__46761;
    wire N__46760;
    wire N__46759;
    wire N__46758;
    wire N__46757;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46739;
    wire N__46736;
    wire N__46733;
    wire N__46730;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46718;
    wire N__46713;
    wire N__46710;
    wire N__46705;
    wire N__46700;
    wire N__46691;
    wire N__46690;
    wire N__46689;
    wire N__46688;
    wire N__46687;
    wire N__46686;
    wire N__46685;
    wire N__46684;
    wire N__46681;
    wire N__46678;
    wire N__46669;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46610;
    wire N__46601;
    wire N__46592;
    wire N__46587;
    wire N__46586;
    wire N__46585;
    wire N__46584;
    wire N__46583;
    wire N__46582;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46578;
    wire N__46577;
    wire N__46576;
    wire N__46573;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46538;
    wire N__46535;
    wire N__46526;
    wire N__46517;
    wire N__46510;
    wire N__46501;
    wire N__46494;
    wire N__46491;
    wire N__46490;
    wire N__46489;
    wire N__46488;
    wire N__46487;
    wire N__46486;
    wire N__46485;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46481;
    wire N__46480;
    wire N__46479;
    wire N__46478;
    wire N__46475;
    wire N__46468;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46446;
    wire N__46445;
    wire N__46444;
    wire N__46443;
    wire N__46442;
    wire N__46439;
    wire N__46436;
    wire N__46429;
    wire N__46420;
    wire N__46417;
    wire N__46412;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46394;
    wire N__46393;
    wire N__46390;
    wire N__46389;
    wire N__46386;
    wire N__46385;
    wire N__46382;
    wire N__46381;
    wire N__46380;
    wire N__46377;
    wire N__46376;
    wire N__46373;
    wire N__46372;
    wire N__46369;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46361;
    wire N__46358;
    wire N__46357;
    wire N__46354;
    wire N__46353;
    wire N__46350;
    wire N__46349;
    wire N__46348;
    wire N__46347;
    wire N__46346;
    wire N__46345;
    wire N__46344;
    wire N__46343;
    wire N__46342;
    wire N__46335;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46317;
    wire N__46308;
    wire N__46307;
    wire N__46306;
    wire N__46305;
    wire N__46304;
    wire N__46301;
    wire N__46294;
    wire N__46289;
    wire N__46286;
    wire N__46283;
    wire N__46278;
    wire N__46263;
    wire N__46246;
    wire N__46229;
    wire N__46222;
    wire N__46213;
    wire N__46210;
    wire N__46201;
    wire N__46198;
    wire N__46193;
    wire N__46190;
    wire N__46187;
    wire N__46182;
    wire N__46177;
    wire N__46162;
    wire N__46159;
    wire N__46154;
    wire N__46151;
    wire N__46146;
    wire N__46145;
    wire N__46144;
    wire N__46143;
    wire N__46142;
    wire N__46139;
    wire N__46134;
    wire N__46125;
    wire N__46122;
    wire N__46117;
    wire N__46114;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46073;
    wire N__46070;
    wire N__46067;
    wire N__46064;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46052;
    wire N__46049;
    wire N__46046;
    wire N__46041;
    wire N__46038;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46026;
    wire N__46023;
    wire N__46022;
    wire N__46019;
    wire N__46016;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45953;
    wire N__45950;
    wire N__45947;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45924;
    wire N__45921;
    wire N__45918;
    wire N__45915;
    wire N__45914;
    wire N__45911;
    wire N__45908;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45885;
    wire N__45882;
    wire N__45881;
    wire N__45878;
    wire N__45875;
    wire N__45870;
    wire N__45867;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45855;
    wire N__45852;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45788;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45764;
    wire N__45761;
    wire N__45758;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45726;
    wire N__45723;
    wire N__45722;
    wire N__45719;
    wire N__45716;
    wire N__45713;
    wire N__45710;
    wire N__45705;
    wire N__45702;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45660;
    wire N__45657;
    wire N__45654;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45483;
    wire N__45480;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45444;
    wire N__45441;
    wire N__45440;
    wire N__45439;
    wire N__45438;
    wire N__45435;
    wire N__45434;
    wire N__45431;
    wire N__45430;
    wire N__45427;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45407;
    wire N__45406;
    wire N__45401;
    wire N__45398;
    wire N__45395;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45351;
    wire N__45348;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45026;
    wire N__45023;
    wire N__45020;
    wire N__45015;
    wire N__45012;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44996;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44973;
    wire N__44972;
    wire N__44971;
    wire N__44970;
    wire N__44969;
    wire N__44968;
    wire N__44967;
    wire N__44966;
    wire N__44965;
    wire N__44964;
    wire N__44963;
    wire N__44962;
    wire N__44961;
    wire N__44960;
    wire N__44959;
    wire N__44958;
    wire N__44957;
    wire N__44956;
    wire N__44955;
    wire N__44954;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44944;
    wire N__44937;
    wire N__44920;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44894;
    wire N__44889;
    wire N__44882;
    wire N__44879;
    wire N__44876;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44852;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44814;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44759;
    wire N__44758;
    wire N__44757;
    wire N__44756;
    wire N__44755;
    wire N__44754;
    wire N__44753;
    wire N__44752;
    wire N__44751;
    wire N__44742;
    wire N__44733;
    wire N__44728;
    wire N__44723;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44711;
    wire N__44708;
    wire N__44705;
    wire N__44700;
    wire N__44699;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44687;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44669;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44648;
    wire N__44645;
    wire N__44642;
    wire N__44637;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44577;
    wire N__44576;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44564;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44528;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44486;
    wire N__44481;
    wire N__44478;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44437;
    wire N__44432;
    wire N__44429;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44419;
    wire N__44414;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44391;
    wire N__44388;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44335;
    wire N__44332;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44306;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44280;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44268;
    wire N__44265;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44241;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44229;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44192;
    wire N__44189;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44157;
    wire N__44154;
    wire N__44153;
    wire N__44150;
    wire N__44147;
    wire N__44144;
    wire N__44141;
    wire N__44138;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44112;
    wire N__44111;
    wire N__44110;
    wire N__44109;
    wire N__44108;
    wire N__44107;
    wire N__44106;
    wire N__44105;
    wire N__44104;
    wire N__44103;
    wire N__44102;
    wire N__44101;
    wire N__44100;
    wire N__44099;
    wire N__44098;
    wire N__44097;
    wire N__44096;
    wire N__44095;
    wire N__44094;
    wire N__44093;
    wire N__44092;
    wire N__44087;
    wire N__44078;
    wire N__44075;
    wire N__44074;
    wire N__44073;
    wire N__44072;
    wire N__44071;
    wire N__44070;
    wire N__44069;
    wire N__44066;
    wire N__44061;
    wire N__44054;
    wire N__44051;
    wire N__44048;
    wire N__44045;
    wire N__44044;
    wire N__44043;
    wire N__44042;
    wire N__44037;
    wire N__44030;
    wire N__44023;
    wire N__44020;
    wire N__44009;
    wire N__44002;
    wire N__43995;
    wire N__43990;
    wire N__43987;
    wire N__43968;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43953;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43932;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43827;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43800;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43785;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43733;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43703;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43686;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43664;
    wire N__43659;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43590;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43574;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43559;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43538;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43526;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43485;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43470;
    wire N__43469;
    wire N__43468;
    wire N__43467;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43435;
    wire N__43432;
    wire N__43425;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43313;
    wire N__43310;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43191;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43155;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43125;
    wire N__43122;
    wire N__43121;
    wire N__43118;
    wire N__43115;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43089;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43002;
    wire N__42999;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42963;
    wire N__42960;
    wire N__42957;
    wire N__42954;
    wire N__42951;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42939;
    wire N__42936;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42798;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42779;
    wire N__42776;
    wire N__42773;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42662;
    wire N__42659;
    wire N__42656;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42575;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42504;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42413;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42403;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42378;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42314;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42296;
    wire N__42295;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42281;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42268;
    wire N__42265;
    wire N__42262;
    wire N__42257;
    wire N__42254;
    wire N__42249;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42223;
    wire N__42220;
    wire N__42217;
    wire N__42214;
    wire N__42207;
    wire N__42206;
    wire N__42201;
    wire N__42198;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42186;
    wire N__42183;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42175;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42159;
    wire N__42158;
    wire N__42157;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42147;
    wire N__42144;
    wire N__42139;
    wire N__42136;
    wire N__42135;
    wire N__42128;
    wire N__42125;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42113;
    wire N__42108;
    wire N__42105;
    wire N__42104;
    wire N__42101;
    wire N__42098;
    wire N__42093;
    wire N__42092;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42005;
    wire N__42002;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41846;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41831;
    wire N__41826;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41811;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41799;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41789;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41774;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41759;
    wire N__41754;
    wire N__41751;
    wire N__41750;
    wire N__41745;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41730;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41718;
    wire N__41717;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41684;
    wire N__41679;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41669;
    wire N__41664;
    wire N__41663;
    wire N__41658;
    wire N__41655;
    wire N__41654;
    wire N__41651;
    wire N__41648;
    wire N__41643;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41605;
    wire N__41602;
    wire N__41599;
    wire N__41596;
    wire N__41593;
    wire N__41590;
    wire N__41583;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41565;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41550;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41522;
    wire N__41517;
    wire N__41514;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41502;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41487;
    wire N__41486;
    wire N__41481;
    wire N__41480;
    wire N__41477;
    wire N__41474;
    wire N__41471;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41441;
    wire N__41436;
    wire N__41433;
    wire N__41432;
    wire N__41427;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41412;
    wire N__41411;
    wire N__41408;
    wire N__41405;
    wire N__41400;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41352;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41330;
    wire N__41325;
    wire N__41322;
    wire N__41321;
    wire N__41316;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41301;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41289;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41267;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41243;
    wire N__41242;
    wire N__41239;
    wire N__41234;
    wire N__41229;
    wire N__41228;
    wire N__41227;
    wire N__41224;
    wire N__41219;
    wire N__41218;
    wire N__41217;
    wire N__41212;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41182;
    wire N__41179;
    wire N__41172;
    wire N__41171;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41156;
    wire N__41153;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41069;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41028;
    wire N__41025;
    wire N__41024;
    wire N__41023;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41007;
    wire N__41004;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40992;
    wire N__40989;
    wire N__40988;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40971;
    wire N__40968;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40956;
    wire N__40955;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40940;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40893;
    wire N__40892;
    wire N__40891;
    wire N__40888;
    wire N__40887;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40869;
    wire N__40866;
    wire N__40865;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40841;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40817;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40800;
    wire N__40797;
    wire N__40796;
    wire N__40795;
    wire N__40792;
    wire N__40787;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40775;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40758;
    wire N__40755;
    wire N__40754;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40739;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40727;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40679;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40662;
    wire N__40659;
    wire N__40656;
    wire N__40655;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40638;
    wire N__40635;
    wire N__40634;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40593;
    wire N__40590;
    wire N__40589;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40574;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40562;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40538;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40514;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40504;
    wire N__40497;
    wire N__40494;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40446;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40438;
    wire N__40433;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40421;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40411;
    wire N__40404;
    wire N__40401;
    wire N__40400;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40390;
    wire N__40385;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40373;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40349;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40339;
    wire N__40332;
    wire N__40329;
    wire N__40328;
    wire N__40325;
    wire N__40322;
    wire N__40317;
    wire N__40314;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40302;
    wire N__40299;
    wire N__40298;
    wire N__40295;
    wire N__40292;
    wire N__40287;
    wire N__40284;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40266;
    wire N__40263;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40244;
    wire N__40241;
    wire N__40238;
    wire N__40233;
    wire N__40230;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40218;
    wire N__40215;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40203;
    wire N__40200;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40188;
    wire N__40185;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40173;
    wire N__40170;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40158;
    wire N__40155;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40143;
    wire N__40140;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40122;
    wire N__40119;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40068;
    wire N__40065;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40053;
    wire N__40050;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40038;
    wire N__40035;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40023;
    wire N__40020;
    wire N__40019;
    wire N__40016;
    wire N__40013;
    wire N__40008;
    wire N__40005;
    wire N__40004;
    wire N__40001;
    wire N__39998;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39960;
    wire N__39957;
    wire N__39956;
    wire N__39953;
    wire N__39950;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39927;
    wire N__39924;
    wire N__39923;
    wire N__39920;
    wire N__39917;
    wire N__39912;
    wire N__39909;
    wire N__39908;
    wire N__39903;
    wire N__39902;
    wire N__39899;
    wire N__39896;
    wire N__39893;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39881;
    wire N__39876;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39861;
    wire N__39858;
    wire N__39857;
    wire N__39854;
    wire N__39851;
    wire N__39850;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39834;
    wire N__39831;
    wire N__39830;
    wire N__39829;
    wire N__39828;
    wire N__39827;
    wire N__39826;
    wire N__39825;
    wire N__39824;
    wire N__39823;
    wire N__39822;
    wire N__39821;
    wire N__39820;
    wire N__39819;
    wire N__39818;
    wire N__39817;
    wire N__39816;
    wire N__39815;
    wire N__39814;
    wire N__39813;
    wire N__39812;
    wire N__39811;
    wire N__39810;
    wire N__39809;
    wire N__39808;
    wire N__39807;
    wire N__39806;
    wire N__39805;
    wire N__39804;
    wire N__39803;
    wire N__39802;
    wire N__39801;
    wire N__39800;
    wire N__39791;
    wire N__39782;
    wire N__39773;
    wire N__39764;
    wire N__39755;
    wire N__39746;
    wire N__39737;
    wire N__39728;
    wire N__39723;
    wire N__39708;
    wire N__39705;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39697;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39681;
    wire N__39680;
    wire N__39679;
    wire N__39676;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39649;
    wire N__39646;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39590;
    wire N__39587;
    wire N__39582;
    wire N__39579;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39542;
    wire N__39541;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39525;
    wire N__39522;
    wire N__39521;
    wire N__39516;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39501;
    wire N__39498;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39483;
    wire N__39480;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39444;
    wire N__39441;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39426;
    wire N__39423;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39408;
    wire N__39405;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39363;
    wire N__39360;
    wire N__39359;
    wire N__39356;
    wire N__39353;
    wire N__39350;
    wire N__39345;
    wire N__39342;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39332;
    wire N__39327;
    wire N__39324;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39309;
    wire N__39306;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39291;
    wire N__39288;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39273;
    wire N__39270;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39255;
    wire N__39252;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39230;
    wire N__39227;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39209;
    wire N__39208;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39197;
    wire N__39194;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39176;
    wire N__39173;
    wire N__39168;
    wire N__39159;
    wire N__39158;
    wire N__39157;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39145;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39092;
    wire N__39087;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39072;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38929;
    wire N__38924;
    wire N__38919;
    wire N__38918;
    wire N__38915;
    wire N__38914;
    wire N__38913;
    wire N__38908;
    wire N__38903;
    wire N__38898;
    wire N__38897;
    wire N__38896;
    wire N__38893;
    wire N__38888;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38771;
    wire N__38766;
    wire N__38763;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38567;
    wire N__38564;
    wire N__38561;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38549;
    wire N__38546;
    wire N__38543;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38424;
    wire N__38423;
    wire N__38420;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38409;
    wire N__38406;
    wire N__38405;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38375;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38342;
    wire N__38341;
    wire N__38338;
    wire N__38333;
    wire N__38328;
    wire N__38327;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38312;
    wire N__38309;
    wire N__38304;
    wire N__38301;
    wire N__38300;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38288;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38261;
    wire N__38260;
    wire N__38257;
    wire N__38252;
    wire N__38247;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38219;
    wire N__38216;
    wire N__38215;
    wire N__38214;
    wire N__38213;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38169;
    wire N__38166;
    wire N__38165;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38151;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38132;
    wire N__38129;
    wire N__38126;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38090;
    wire N__38089;
    wire N__38088;
    wire N__38087;
    wire N__38086;
    wire N__38085;
    wire N__38084;
    wire N__38083;
    wire N__38082;
    wire N__38081;
    wire N__38080;
    wire N__38079;
    wire N__38078;
    wire N__38077;
    wire N__38076;
    wire N__38075;
    wire N__38074;
    wire N__38073;
    wire N__38072;
    wire N__38067;
    wire N__38058;
    wire N__38057;
    wire N__38056;
    wire N__38055;
    wire N__38054;
    wire N__38045;
    wire N__38036;
    wire N__38027;
    wire N__38018;
    wire N__38009;
    wire N__38004;
    wire N__37995;
    wire N__37982;
    wire N__37977;
    wire N__37974;
    wire N__37973;
    wire N__37972;
    wire N__37969;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37951;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37922;
    wire N__37921;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37905;
    wire N__37904;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37868;
    wire N__37867;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37739;
    wire N__37738;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37720;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37356;
    wire N__37353;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37266;
    wire N__37263;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37155;
    wire N__37152;
    wire N__37149;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37106;
    wire N__37103;
    wire N__37102;
    wire N__37095;
    wire N__37092;
    wire N__37091;
    wire N__37086;
    wire N__37083;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37072;
    wire N__37067;
    wire N__37064;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37040;
    wire N__37037;
    wire N__37036;
    wire N__37033;
    wire N__37032;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37017;
    wire N__37014;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36985;
    wire N__36978;
    wire N__36975;
    wire N__36974;
    wire N__36971;
    wire N__36970;
    wire N__36967;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36921;
    wire N__36912;
    wire N__36911;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36885;
    wire N__36882;
    wire N__36881;
    wire N__36878;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36866;
    wire N__36863;
    wire N__36858;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36846;
    wire N__36845;
    wire N__36844;
    wire N__36843;
    wire N__36840;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36822;
    wire N__36821;
    wire N__36818;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36787;
    wire N__36784;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36759;
    wire N__36758;
    wire N__36755;
    wire N__36754;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36739;
    wire N__36736;
    wire N__36729;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36708;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36681;
    wire N__36678;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36657;
    wire N__36654;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36646;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36615;
    wire N__36612;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36590;
    wire N__36589;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36567;
    wire N__36566;
    wire N__36565;
    wire N__36562;
    wire N__36557;
    wire N__36550;
    wire N__36547;
    wire N__36542;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36530;
    wire N__36529;
    wire N__36526;
    wire N__36521;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36505;
    wire N__36502;
    wire N__36497;
    wire N__36494;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36462;
    wire N__36461;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36414;
    wire N__36411;
    wire N__36408;
    wire N__36407;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36392;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36377;
    wire N__36374;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36335;
    wire N__36334;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36314;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36276;
    wire N__36271;
    wire N__36266;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36248;
    wire N__36247;
    wire N__36244;
    wire N__36239;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36223;
    wire N__36222;
    wire N__36221;
    wire N__36214;
    wire N__36213;
    wire N__36212;
    wire N__36211;
    wire N__36210;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36205;
    wire N__36204;
    wire N__36203;
    wire N__36202;
    wire N__36201;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36184;
    wire N__36175;
    wire N__36172;
    wire N__36163;
    wire N__36154;
    wire N__36145;
    wire N__36134;
    wire N__36125;
    wire N__36114;
    wire N__36109;
    wire N__36102;
    wire N__36099;
    wire N__36098;
    wire N__36097;
    wire N__36094;
    wire N__36089;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36077;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36062;
    wire N__36059;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36042;
    wire N__36041;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35939;
    wire N__35938;
    wire N__35935;
    wire N__35930;
    wire N__35925;
    wire N__35922;
    wire N__35921;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35904;
    wire N__35901;
    wire N__35900;
    wire N__35897;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35887;
    wire N__35880;
    wire N__35877;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35863;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35840;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35810;
    wire N__35807;
    wire N__35806;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35790;
    wire N__35787;
    wire N__35786;
    wire N__35783;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35760;
    wire N__35757;
    wire N__35756;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35739;
    wire N__35736;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35732;
    wire N__35731;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35727;
    wire N__35726;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35722;
    wire N__35721;
    wire N__35720;
    wire N__35719;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35709;
    wire N__35708;
    wire N__35707;
    wire N__35706;
    wire N__35705;
    wire N__35696;
    wire N__35689;
    wire N__35680;
    wire N__35669;
    wire N__35660;
    wire N__35651;
    wire N__35642;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35616;
    wire N__35613;
    wire N__35606;
    wire N__35601;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35577;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35531;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35514;
    wire N__35511;
    wire N__35510;
    wire N__35507;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35490;
    wire N__35487;
    wire N__35486;
    wire N__35485;
    wire N__35482;
    wire N__35477;
    wire N__35472;
    wire N__35469;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35454;
    wire N__35451;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35436;
    wire N__35433;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35415;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35382;
    wire N__35379;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35364;
    wire N__35361;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35346;
    wire N__35343;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35328;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35286;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35247;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35232;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35175;
    wire N__35172;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35136;
    wire N__35133;
    wire N__35132;
    wire N__35129;
    wire N__35126;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35114;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34908;
    wire N__34907;
    wire N__34906;
    wire N__34905;
    wire N__34904;
    wire N__34903;
    wire N__34902;
    wire N__34901;
    wire N__34900;
    wire N__34899;
    wire N__34898;
    wire N__34897;
    wire N__34894;
    wire N__34893;
    wire N__34888;
    wire N__34887;
    wire N__34884;
    wire N__34871;
    wire N__34866;
    wire N__34861;
    wire N__34860;
    wire N__34859;
    wire N__34858;
    wire N__34857;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34850;
    wire N__34849;
    wire N__34848;
    wire N__34847;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34840;
    wire N__34835;
    wire N__34832;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34811;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34794;
    wire N__34793;
    wire N__34792;
    wire N__34791;
    wire N__34788;
    wire N__34787;
    wire N__34786;
    wire N__34785;
    wire N__34784;
    wire N__34783;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34775;
    wire N__34774;
    wire N__34773;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34763;
    wire N__34762;
    wire N__34759;
    wire N__34758;
    wire N__34755;
    wire N__34754;
    wire N__34751;
    wire N__34750;
    wire N__34747;
    wire N__34746;
    wire N__34745;
    wire N__34744;
    wire N__34743;
    wire N__34742;
    wire N__34741;
    wire N__34740;
    wire N__34739;
    wire N__34738;
    wire N__34737;
    wire N__34736;
    wire N__34735;
    wire N__34734;
    wire N__34733;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34712;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34686;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34678;
    wire N__34677;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34647;
    wire N__34644;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34640;
    wire N__34639;
    wire N__34638;
    wire N__34637;
    wire N__34630;
    wire N__34625;
    wire N__34622;
    wire N__34621;
    wire N__34618;
    wire N__34617;
    wire N__34614;
    wire N__34613;
    wire N__34596;
    wire N__34593;
    wire N__34592;
    wire N__34589;
    wire N__34588;
    wire N__34585;
    wire N__34584;
    wire N__34581;
    wire N__34580;
    wire N__34577;
    wire N__34576;
    wire N__34573;
    wire N__34572;
    wire N__34569;
    wire N__34568;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34560;
    wire N__34559;
    wire N__34556;
    wire N__34555;
    wire N__34552;
    wire N__34551;
    wire N__34550;
    wire N__34547;
    wire N__34546;
    wire N__34543;
    wire N__34542;
    wire N__34539;
    wire N__34538;
    wire N__34529;
    wire N__34526;
    wire N__34517;
    wire N__34508;
    wire N__34505;
    wire N__34494;
    wire N__34493;
    wire N__34492;
    wire N__34491;
    wire N__34490;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34474;
    wire N__34471;
    wire N__34470;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34462;
    wire N__34459;
    wire N__34458;
    wire N__34455;
    wire N__34454;
    wire N__34451;
    wire N__34450;
    wire N__34447;
    wire N__34446;
    wire N__34441;
    wire N__34428;
    wire N__34425;
    wire N__34408;
    wire N__34391;
    wire N__34376;
    wire N__34373;
    wire N__34360;
    wire N__34357;
    wire N__34346;
    wire N__34337;
    wire N__34328;
    wire N__34311;
    wire N__34298;
    wire N__34281;
    wire N__34266;
    wire N__34265;
    wire N__34264;
    wire N__34261;
    wire N__34260;
    wire N__34259;
    wire N__34258;
    wire N__34255;
    wire N__34254;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34242;
    wire N__34239;
    wire N__34238;
    wire N__34237;
    wire N__34236;
    wire N__34235;
    wire N__34234;
    wire N__34231;
    wire N__34230;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34215;
    wire N__34212;
    wire N__34211;
    wire N__34210;
    wire N__34209;
    wire N__34208;
    wire N__34203;
    wire N__34202;
    wire N__34201;
    wire N__34200;
    wire N__34199;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34188;
    wire N__34187;
    wire N__34186;
    wire N__34185;
    wire N__34182;
    wire N__34177;
    wire N__34174;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34153;
    wire N__34148;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34136;
    wire N__34135;
    wire N__34134;
    wire N__34133;
    wire N__34130;
    wire N__34117;
    wire N__34100;
    wire N__34091;
    wire N__34090;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34079;
    wire N__34078;
    wire N__34077;
    wire N__34076;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34072;
    wire N__34071;
    wire N__34070;
    wire N__34069;
    wire N__34068;
    wire N__34067;
    wire N__34066;
    wire N__34065;
    wire N__34064;
    wire N__34063;
    wire N__34062;
    wire N__34061;
    wire N__34060;
    wire N__34057;
    wire N__34046;
    wire N__34039;
    wire N__34034;
    wire N__34027;
    wire N__34018;
    wire N__34015;
    wire N__34006;
    wire N__34001;
    wire N__33998;
    wire N__33985;
    wire N__33974;
    wire N__33961;
    wire N__33956;
    wire N__33949;
    wire N__33942;
    wire N__33921;
    wire N__33918;
    wire N__33917;
    wire N__33916;
    wire N__33915;
    wire N__33912;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33887;
    wire N__33882;
    wire N__33881;
    wire N__33880;
    wire N__33877;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33776;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33758;
    wire N__33757;
    wire N__33756;
    wire N__33755;
    wire N__33754;
    wire N__33753;
    wire N__33752;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33652;
    wire N__33647;
    wire N__33642;
    wire N__33639;
    wire N__33638;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33589;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33545;
    wire N__33544;
    wire N__33541;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33513;
    wire N__33510;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33439;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33416;
    wire N__33411;
    wire N__33410;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33357;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33338;
    wire N__33333;
    wire N__33332;
    wire N__33329;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33212;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33185;
    wire N__33182;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33162;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33140;
    wire N__33137;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33104;
    wire N__33101;
    wire N__33100;
    wire N__33097;
    wire N__33096;
    wire N__33095;
    wire N__33094;
    wire N__33091;
    wire N__33086;
    wire N__33083;
    wire N__33078;
    wire N__33075;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32972;
    wire N__32971;
    wire N__32968;
    wire N__32963;
    wire N__32958;
    wire N__32955;
    wire N__32954;
    wire N__32953;
    wire N__32950;
    wire N__32945;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32897;
    wire N__32892;
    wire N__32889;
    wire N__32888;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32876;
    wire N__32873;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32850;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32822;
    wire N__32817;
    wire N__32816;
    wire N__32815;
    wire N__32810;
    wire N__32807;
    wire N__32802;
    wire N__32801;
    wire N__32800;
    wire N__32799;
    wire N__32798;
    wire N__32797;
    wire N__32794;
    wire N__32789;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32761;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32697;
    wire N__32696;
    wire N__32695;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32557;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32328;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32277;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32252;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32235;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32197;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32182;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32150;
    wire N__32149;
    wire N__32146;
    wire N__32141;
    wire N__32140;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32102;
    wire N__32099;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32088;
    wire N__32085;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32069;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32013;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31958;
    wire N__31955;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31939;
    wire N__31936;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31886;
    wire N__31883;
    wire N__31882;
    wire N__31879;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31858;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31826;
    wire N__31825;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31795;
    wire N__31792;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31757;
    wire N__31756;
    wire N__31753;
    wire N__31748;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31690;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31669;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31655;
    wire N__31654;
    wire N__31653;
    wire N__31652;
    wire N__31651;
    wire N__31650;
    wire N__31649;
    wire N__31648;
    wire N__31647;
    wire N__31644;
    wire N__31643;
    wire N__31642;
    wire N__31641;
    wire N__31640;
    wire N__31637;
    wire N__31636;
    wire N__31635;
    wire N__31626;
    wire N__31617;
    wire N__31614;
    wire N__31613;
    wire N__31610;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31594;
    wire N__31593;
    wire N__31592;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31588;
    wire N__31587;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31582;
    wire N__31579;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31563;
    wire N__31560;
    wire N__31555;
    wire N__31552;
    wire N__31545;
    wire N__31542;
    wire N__31535;
    wire N__31522;
    wire N__31517;
    wire N__31514;
    wire N__31505;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31420;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31399;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31361;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31350;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31307;
    wire N__31304;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31267;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31193;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31157;
    wire N__31156;
    wire N__31155;
    wire N__31152;
    wire N__31147;
    wire N__31144;
    wire N__31139;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31115;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31084;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31042;
    wire N__31041;
    wire N__31038;
    wire N__31033;
    wire N__31030;
    wire N__31025;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30978;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30835;
    wire N__30830;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30794;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30774;
    wire N__30771;
    wire N__30766;
    wire N__30763;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30731;
    wire N__30728;
    wire N__30727;
    wire N__30724;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30694;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30656;
    wire N__30655;
    wire N__30652;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30548;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30508;
    wire N__30505;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30482;
    wire N__30479;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30445;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30431;
    wire N__30428;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30352;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30334;
    wire N__30331;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30295;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30232;
    wire N__30229;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30173;
    wire N__30172;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30106;
    wire N__30105;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30059;
    wire N__30058;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30023;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30008;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29971;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29945;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29930;
    wire N__29925;
    wire N__29922;
    wire N__29921;
    wire N__29918;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29900;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29881;
    wire N__29880;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29865;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29849;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29822;
    wire N__29819;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29771;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29717;
    wire N__29714;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29672;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29636;
    wire N__29633;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29594;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29429;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29386;
    wire N__29381;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29357;
    wire N__29356;
    wire N__29353;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29310;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29189;
    wire N__29186;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29114;
    wire N__29113;
    wire N__29110;
    wire N__29105;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29087;
    wire N__29084;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29066;
    wire N__29061;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29042;
    wire N__29041;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28967;
    wire N__28962;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28953;
    wire N__28952;
    wire N__28951;
    wire N__28950;
    wire N__28949;
    wire N__28948;
    wire N__28947;
    wire N__28946;
    wire N__28945;
    wire N__28944;
    wire N__28943;
    wire N__28940;
    wire N__28931;
    wire N__28924;
    wire N__28911;
    wire N__28910;
    wire N__28909;
    wire N__28908;
    wire N__28901;
    wire N__28894;
    wire N__28891;
    wire N__28884;
    wire N__28883;
    wire N__28882;
    wire N__28881;
    wire N__28880;
    wire N__28877;
    wire N__28876;
    wire N__28873;
    wire N__28868;
    wire N__28863;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28832;
    wire N__28829;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28802;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28789;
    wire N__28782;
    wire N__28779;
    wire N__28778;
    wire N__28777;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28766;
    wire N__28765;
    wire N__28762;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28740;
    wire N__28731;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28704;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28680;
    wire N__28679;
    wire N__28678;
    wire N__28675;
    wire N__28670;
    wire N__28665;
    wire N__28664;
    wire N__28663;
    wire N__28660;
    wire N__28655;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28631;
    wire N__28630;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28614;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28606;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28559;
    wire N__28558;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28542;
    wire N__28541;
    wire N__28540;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28469;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28452;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28418;
    wire N__28417;
    wire N__28416;
    wire N__28413;
    wire N__28408;
    wire N__28405;
    wire N__28398;
    wire N__28397;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28380;
    wire N__28379;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28061;
    wire N__28056;
    wire N__28055;
    wire N__28052;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28035;
    wire N__28034;
    wire N__28033;
    wire N__28030;
    wire N__28029;
    wire N__28028;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__27999;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27969;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27905;
    wire N__27902;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27885;
    wire N__27882;
    wire N__27881;
    wire N__27878;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27854;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27837;
    wire N__27834;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27822;
    wire N__27821;
    wire N__27818;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27801;
    wire N__27798;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27786;
    wire N__27785;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27758;
    wire N__27755;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27738;
    wire N__27735;
    wire N__27734;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27723;
    wire N__27718;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27702;
    wire N__27699;
    wire N__27698;
    wire N__27695;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27678;
    wire N__27677;
    wire N__27674;
    wire N__27673;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27641;
    wire N__27636;
    wire N__27633;
    wire N__27632;
    wire N__27629;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27612;
    wire N__27609;
    wire N__27608;
    wire N__27605;
    wire N__27604;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27570;
    wire N__27567;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27546;
    wire N__27545;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27523;
    wire N__27518;
    wire N__27513;
    wire N__27510;
    wire N__27509;
    wire N__27506;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27474;
    wire N__27471;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27455;
    wire N__27450;
    wire N__27447;
    wire N__27446;
    wire N__27443;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27426;
    wire N__27423;
    wire N__27422;
    wire N__27419;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27402;
    wire N__27399;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27378;
    wire N__27375;
    wire N__27374;
    wire N__27371;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27354;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27330;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27318;
    wire N__27315;
    wire N__27314;
    wire N__27311;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27257;
    wire N__27252;
    wire N__27249;
    wire N__27248;
    wire N__27245;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27228;
    wire N__27227;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27190;
    wire N__27183;
    wire N__27180;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27159;
    wire N__27156;
    wire N__27155;
    wire N__27152;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27135;
    wire N__27132;
    wire N__27131;
    wire N__27128;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27111;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27103;
    wire N__27100;
    wire N__27095;
    wire N__27094;
    wire N__27089;
    wire N__27086;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27074;
    wire N__27071;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27054;
    wire N__27051;
    wire N__27050;
    wire N__27047;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26983;
    wire N__26976;
    wire N__26973;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26965;
    wire N__26964;
    wire N__26959;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26943;
    wire N__26940;
    wire N__26939;
    wire N__26936;
    wire N__26935;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26894;
    wire N__26889;
    wire N__26886;
    wire N__26885;
    wire N__26882;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26865;
    wire N__26862;
    wire N__26861;
    wire N__26858;
    wire N__26857;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26834;
    wire N__26829;
    wire N__26826;
    wire N__26825;
    wire N__26822;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26805;
    wire N__26804;
    wire N__26803;
    wire N__26800;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26771;
    wire N__26768;
    wire N__26763;
    wire N__26760;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26734;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26713;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26696;
    wire N__26693;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26294;
    wire N__26293;
    wire N__26292;
    wire N__26291;
    wire N__26290;
    wire N__26289;
    wire N__26288;
    wire N__26287;
    wire N__26286;
    wire N__26285;
    wire N__26284;
    wire N__26283;
    wire N__26282;
    wire N__26281;
    wire N__26280;
    wire N__26279;
    wire N__26278;
    wire N__26277;
    wire N__26276;
    wire N__26275;
    wire N__26274;
    wire N__26273;
    wire N__26272;
    wire N__26271;
    wire N__26270;
    wire N__26269;
    wire N__26268;
    wire N__26267;
    wire N__26266;
    wire N__26265;
    wire N__26264;
    wire N__26255;
    wire N__26246;
    wire N__26237;
    wire N__26228;
    wire N__26219;
    wire N__26210;
    wire N__26201;
    wire N__26192;
    wire N__26183;
    wire N__26172;
    wire N__26169;
    wire N__26168;
    wire N__26167;
    wire N__26166;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26121;
    wire N__26118;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26106;
    wire N__26103;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25973;
    wire N__25972;
    wire N__25971;
    wire N__25970;
    wire N__25969;
    wire N__25968;
    wire N__25967;
    wire N__25966;
    wire N__25965;
    wire N__25964;
    wire N__25963;
    wire N__25962;
    wire N__25961;
    wire N__25960;
    wire N__25959;
    wire N__25958;
    wire N__25957;
    wire N__25956;
    wire N__25955;
    wire N__25954;
    wire N__25953;
    wire N__25948;
    wire N__25947;
    wire N__25946;
    wire N__25945;
    wire N__25944;
    wire N__25935;
    wire N__25934;
    wire N__25933;
    wire N__25932;
    wire N__25931;
    wire N__25922;
    wire N__25913;
    wire N__25904;
    wire N__25895;
    wire N__25892;
    wire N__25883;
    wire N__25880;
    wire N__25871;
    wire N__25862;
    wire N__25857;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25841;
    wire N__25840;
    wire N__25837;
    wire N__25832;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25801;
    wire N__25798;
    wire N__25797;
    wire N__25790;
    wire N__25787;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25661;
    wire N__25658;
    wire N__25657;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25273;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25241;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25213;
    wire N__25208;
    wire N__25205;
    wire N__25200;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24593;
    wire N__24592;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24586;
    wire N__24585;
    wire N__24584;
    wire N__24583;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24579;
    wire N__24574;
    wire N__24569;
    wire N__24566;
    wire N__24565;
    wire N__24564;
    wire N__24563;
    wire N__24562;
    wire N__24561;
    wire N__24560;
    wire N__24559;
    wire N__24558;
    wire N__24555;
    wire N__24544;
    wire N__24541;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24535;
    wire N__24534;
    wire N__24533;
    wire N__24528;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24501;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24483;
    wire N__24476;
    wire N__24475;
    wire N__24466;
    wire N__24459;
    wire N__24458;
    wire N__24457;
    wire N__24456;
    wire N__24455;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24443;
    wire N__24432;
    wire N__24429;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24071;
    wire N__24070;
    wire N__24063;
    wire N__24060;
    wire N__24059;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23961;
    wire N__23958;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23950;
    wire N__23947;
    wire N__23942;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23886;
    wire N__23883;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23838;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23778;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23490;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23463;
    wire N__23460;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23439;
    wire N__23436;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23379;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23358;
    wire N__23355;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23298;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23280;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23259;
    wire N__23256;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23235;
    wire N__23232;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23211;
    wire N__23208;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23187;
    wire N__23184;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22656;
    wire N__22653;
    wire N__22652;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22647;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22633;
    wire N__22632;
    wire N__22629;
    wire N__22628;
    wire N__22627;
    wire N__22626;
    wire N__22625;
    wire N__22624;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22598;
    wire N__22597;
    wire N__22596;
    wire N__22595;
    wire N__22592;
    wire N__22587;
    wire N__22580;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22559;
    wire N__22558;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22554;
    wire N__22553;
    wire N__22552;
    wire N__22551;
    wire N__22550;
    wire N__22545;
    wire N__22542;
    wire N__22533;
    wire N__22528;
    wire N__22523;
    wire N__22520;
    wire N__22511;
    wire N__22502;
    wire N__22499;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21519;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21511;
    wire N__21510;
    wire N__21509;
    wire N__21508;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21459;
    wire N__21450;
    wire N__21447;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire N_94_i_i;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire bfn_2_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire bfn_2_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire bfn_2_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_2_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire un8_start_stop;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire bfn_3_11_0_;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire bfn_3_12_0_;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire bfn_3_13_0_;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire bfn_3_14_0_;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.N_1571_i ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_77 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.N_46_21 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \current_shift_inst.PI_CTRL.N_46_16_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.control_input_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_5_11_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_5_12_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_5_13_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_5_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire delay_hc_input_c_g;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_4 ;
    wire \phase_controller_inst2.start_flagZ0 ;
    wire \phase_controller_inst2.state_ns_0_0_1 ;
    wire bfn_8_11_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_8_12_0_;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_8_13_0_;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_8_14_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire s4_phy_c;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_start_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire bfn_9_22_0_;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire s3_phy_c;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire bfn_10_7_0_;
    wire \phase_controller_inst2.stoper_tr.counter_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_7 ;
    wire bfn_10_8_0_;
    wire \phase_controller_inst2.stoper_tr.counter_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_15 ;
    wire bfn_10_9_0_;
    wire \phase_controller_inst2.stoper_tr.counter_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_23 ;
    wire bfn_10_10_0_;
    wire \phase_controller_inst2.stoper_tr.counter_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_i_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_g ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_10_20_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_10_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_10_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_10_23_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_start_0 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_0 ;
    wire bfn_11_7_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_1 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_8 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_9 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_15 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_30 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.counter ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_start_0 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire bfn_11_19_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_11_20_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire bfn_11_21_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire bfn_11_22_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_0 ;
    wire bfn_11_25_0_;
    wire \phase_controller_inst1.stoper_tr.counter_i_1 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_8 ;
    wire bfn_11_26_0_;
    wire \phase_controller_inst1.stoper_tr.counter_i_9 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_15 ;
    wire bfn_11_27_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_30 ;
    wire bfn_11_28_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt24 ;
    wire \current_shift_inst.timer_s1.N_154_i ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt26 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ;
    wire delay_tr_input_c_g;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.timer_s1.N_153_i_g ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.counter ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_0 ;
    wire bfn_12_27_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_8 ;
    wire bfn_12_28_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_15 ;
    wire bfn_12_29_0_;
    wire \phase_controller_inst1.stoper_tr.counter_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_24 ;
    wire bfn_12_30_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_i_0 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_g ;
    wire bfn_13_7_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_7 ;
    wire bfn_13_8_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_15 ;
    wire bfn_13_9_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_23 ;
    wire bfn_13_10_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_i_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire il_max_comp1_c;
    wire start_stop_c;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.state_ns_0_0_1_cascade_ ;
    wire \phase_controller_inst1.start_flagZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_start_0 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ;
    wire bfn_13_19_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_1;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_2;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_3;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_4;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_5;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_6;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_7;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_8;
    wire bfn_13_20_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_9;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_10;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_11;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_12;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_13;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_14;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_15;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_16;
    wire bfn_13_21_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_17;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_18;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_20;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_21;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_22;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_23;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_24;
    wire bfn_13_22_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_25;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_26;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_27;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire bfn_13_23_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_13_24_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_13_25_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_13_26_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_158_i ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_19;
    wire \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt18 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \current_shift_inst.timer_s1.N_153_i ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.counter ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_0 ;
    wire bfn_14_8_0_;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_1 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_8 ;
    wire bfn_14_9_0_;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_9 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_15 ;
    wire bfn_14_10_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_30 ;
    wire bfn_14_11_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_0 ;
    wire bfn_14_12_0_;
    wire \phase_controller_inst1.stoper_hc.counter_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_8 ;
    wire bfn_14_13_0_;
    wire \phase_controller_inst1.stoper_hc.counter_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_15 ;
    wire bfn_14_14_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30 ;
    wire bfn_14_15_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNILK91B_0_9_cascade_;
    wire \phase_controller_inst1.stoper_hc.counter ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_0 ;
    wire bfn_14_16_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_8 ;
    wire bfn_14_17_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_15 ;
    wire bfn_14_18_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_23 ;
    wire bfn_14_19_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_i_0 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ;
    wire bfn_14_20_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ;
    wire bfn_14_21_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ;
    wire bfn_14_22_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ;
    wire bfn_14_23_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_28;
    wire bfn_14_24_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_14_25_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_14_26_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_14_27_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire s1_phy_c;
    wire state_3;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire elapsed_time_ns_1_RNIK63T9_0_8_cascade_;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire elapsed_time_ns_1_RNIU0DN9_0_20_cascade_;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire elapsed_time_ns_1_RNIL73T9_0_9_cascade_;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire elapsed_time_ns_1_RNIU7OBB_0_11_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire elapsed_time_ns_1_RNI68CN9_0_19_cascade_;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire elapsed_time_ns_1_RNIV8OBB_0_12_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire elapsed_time_ns_1_RNIV9PBB_0_21_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIIH91B_0_6_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire elapsed_time_ns_1_RNIJI91B_0_7_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_157_i ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire elapsed_time_ns_1_RNIU8PBB_0_20_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire elapsed_time_ns_1_RNI3DOBB_0_16_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire elapsed_time_ns_1_RNIT6OBB_0_10_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI5FOBB_0_18_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire elapsed_time_ns_1_RNI3EPBB_0_25_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire elapsed_time_ns_1_RNI0BPBB_0_22_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire elapsed_time_ns_1_RNI1CPBB_0_23_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire elapsed_time_ns_1_RNIVAQBB_0_30_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire elapsed_time_ns_1_RNI7IPBB_0_29_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire elapsed_time_ns_1_RNI6GOBB_0_19_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire bfn_15_28_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire bfn_15_29_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_15_30_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire elapsed_time_ns_1_RNI57CN9_0_18_cascade_;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire elapsed_time_ns_1_RNIF13T9_0_3_cascade_;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire elapsed_time_ns_1_RNIJ53T9_0_7_cascade_;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire elapsed_time_ns_1_RNI35CN9_0_16_cascade_;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire elapsed_time_ns_1_RNIG23T9_0_4_cascade_;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire elapsed_time_ns_1_RNI24CN9_0_15_cascade_;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire elapsed_time_ns_1_RNI13CN9_0_14_cascade_;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire elapsed_time_ns_1_RNIUVBN9_0_11_cascade_;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire elapsed_time_ns_1_RNI2COBB_0_15_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire elapsed_time_ns_1_RNIGF91B_0_4_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire bfn_16_23_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_16_24_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire pwm_duty_input_10;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_16_28_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_16_29_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire bfn_16_30_0_;
    wire GB_BUFFER_red_c_g_THRU_CO;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ;
    wire bfn_17_8_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_1;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_2;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_3;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_4;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_5;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_6;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_7;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_8;
    wire bfn_17_9_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_9;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_10;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_11;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_12;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_13;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_14;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_15;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ;
    wire bfn_17_10_0_;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_20;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_21;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_22;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_23;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ;
    wire CONSTANT_ONE_NET;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ;
    wire bfn_17_12_0_;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ;
    wire bfn_17_13_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ;
    wire bfn_17_14_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ;
    wire bfn_17_15_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_28;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire bfn_17_16_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_17_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire bfn_17_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_17_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire bfn_17_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_17_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_17_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_17_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_156_i ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_17_24_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_17_25_0_;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.un19_threshold_0_axb_0 ;
    wire \pwm_generator_inst.un14_counter_0 ;
    wire bfn_17_26_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_2 ;
    wire \pwm_generator_inst.un14_counter_2 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_3 ;
    wire \pwm_generator_inst.un14_counter_3 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_2 ;
    wire \pwm_generator_inst.un14_counter_4 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_5 ;
    wire \pwm_generator_inst.un14_counter_5 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_7 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_7 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire bfn_17_27_0_;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_0_cry_8 ;
    wire \pwm_generator_inst.un14_counter_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_0_axb_8 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_16;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_18;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_19;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_17;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_27;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_26;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_24;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_25;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire elapsed_time_ns_1_RNIV0CN9_0_12_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire elapsed_time_ns_1_RNI14DN9_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire elapsed_time_ns_1_RNI58DN9_0_27_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire elapsed_time_ns_1_RNI7ADN9_0_29_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_155_i ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_20_25_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_20_26_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un19_threshold_0_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire bfn_20_27_0_;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire pwm_duty_input_0;
    wire \current_shift_inst.PI_CTRL.N_152 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire pwm_duty_input_3;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire pwm_duty_input_9;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire pwm_duty_input_5;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire pwm_duty_input_8;
    wire \current_shift_inst.PI_CTRL.N_150 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire pwm_duty_input_7;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__21981),
            .RESETB(N__45795),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__46145),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__46142),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__23358,N__23235,N__23990,N__23211,N__23406,N__23187,N__23439,N__23807,N__23723,N__23837,N__23490,N__23259,N__23463,N__23379,N__23064,N__26103}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__46144,dangling_wire_45,N__46143}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__46449),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__46442),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__44966,N__44959,N__44964,N__44958,N__44965,N__44957,N__44967,N__44954,N__44960,N__44953,N__44961,N__44955,N__44962,N__44956,N__44963}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__46448,N__46445,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__46443,N__46447,N__46444,N__46446}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__46586),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__46579),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__44968,N__44971,N__44969,N__44972,N__44970,N__52836,N__52701,N__52509,N__52791,N__52743,N__52878,N__51510,N__51633,N__51576,N__51615}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__46585,N__46582,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__46580,N__46584,N__46581,N__46583}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__46305),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__46304),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__23280,N__26082,N__23297,N__26117,N__23319,N__23855,N__23882,N__23088,N__23622,N__26150,N__23777,N__23517,N__23915,N__23741,N__22673}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__46307,dangling_wire_215,N__46306}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__53074),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__53076),
            .DIN(N__53075),
            .DOUT(N__53074),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__53076),
            .PADOUT(N__53075),
            .PADIN(N__53074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__53065),
            .DIN(N__53064),
            .DOUT(N__53063),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__53065),
            .PADOUT(N__53064),
            .PADIN(N__53063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__49554),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__53056),
            .DIN(N__53055),
            .DOUT(N__53054),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__53056),
            .PADOUT(N__53055),
            .PADIN(N__53054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38235),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__53047),
            .DIN(N__53046),
            .DOUT(N__53045),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__53047),
            .PADOUT(N__53046),
            .PADIN(N__53045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__53038),
            .DIN(N__53037),
            .DOUT(N__53036),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__53038),
            .PADOUT(N__53037),
            .PADIN(N__53036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__41250),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__53029),
            .DIN(N__53028),
            .DOUT(N__53027),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__53029),
            .PADOUT(N__53028),
            .PADIN(N__53027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25044),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__53020),
            .DIN(N__53019),
            .DOUT(N__53018),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__53020),
            .PADOUT(N__53019),
            .PADIN(N__53018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__53011),
            .DIN(N__53010),
            .DOUT(N__53009),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__53011),
            .PADOUT(N__53010),
            .PADIN(N__53009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25812),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__53002),
            .DIN(N__53001),
            .DOUT(N__53000),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__53002),
            .PADOUT(N__53001),
            .PADIN(N__53000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__52993),
            .DIN(N__52992),
            .DOUT(N__52991),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__52993),
            .PADOUT(N__52992),
            .PADIN(N__52991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__52984),
            .DIN(N__52983),
            .DOUT(N__52982),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__52984),
            .PADOUT(N__52983),
            .PADIN(N__52982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__52975),
            .DIN(N__52974),
            .DOUT(N__52973),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__52975),
            .PADOUT(N__52974),
            .PADIN(N__52973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__52966),
            .DIN(N__52965),
            .DOUT(N__52964),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__52966),
            .PADOUT(N__52965),
            .PADIN(N__52964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12380 (
            .O(N__52947),
            .I(N__52944));
    LocalMux I__12379 (
            .O(N__52944),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__12378 (
            .O(N__52941),
            .I(N__52936));
    CascadeMux I__12377 (
            .O(N__52940),
            .I(N__52933));
    CascadeMux I__12376 (
            .O(N__52939),
            .I(N__52930));
    LocalMux I__12375 (
            .O(N__52936),
            .I(N__52926));
    InMux I__12374 (
            .O(N__52933),
            .I(N__52921));
    InMux I__12373 (
            .O(N__52930),
            .I(N__52921));
    InMux I__12372 (
            .O(N__52929),
            .I(N__52918));
    Span4Mux_v I__12371 (
            .O(N__52926),
            .I(N__52915));
    LocalMux I__12370 (
            .O(N__52921),
            .I(N__52910));
    LocalMux I__12369 (
            .O(N__52918),
            .I(N__52910));
    Sp12to4 I__12368 (
            .O(N__52915),
            .I(N__52905));
    Span12Mux_v I__12367 (
            .O(N__52910),
            .I(N__52905));
    Span12Mux_h I__12366 (
            .O(N__52905),
            .I(N__52902));
    Odrv12 I__12365 (
            .O(N__52902),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    CascadeMux I__12364 (
            .O(N__52899),
            .I(N__52896));
    InMux I__12363 (
            .O(N__52896),
            .I(N__52892));
    CascadeMux I__12362 (
            .O(N__52895),
            .I(N__52889));
    LocalMux I__12361 (
            .O(N__52892),
            .I(N__52886));
    InMux I__12360 (
            .O(N__52889),
            .I(N__52883));
    Odrv4 I__12359 (
            .O(N__52886),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__12358 (
            .O(N__52883),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__12357 (
            .O(N__52878),
            .I(N__52875));
    LocalMux I__12356 (
            .O(N__52875),
            .I(N__52872));
    Odrv4 I__12355 (
            .O(N__52872),
            .I(pwm_duty_input_4));
    CascadeMux I__12354 (
            .O(N__52869),
            .I(N__52866));
    InMux I__12353 (
            .O(N__52866),
            .I(N__52863));
    LocalMux I__12352 (
            .O(N__52863),
            .I(N__52858));
    InMux I__12351 (
            .O(N__52862),
            .I(N__52853));
    InMux I__12350 (
            .O(N__52861),
            .I(N__52853));
    Span4Mux_v I__12349 (
            .O(N__52858),
            .I(N__52848));
    LocalMux I__12348 (
            .O(N__52853),
            .I(N__52848));
    Span4Mux_h I__12347 (
            .O(N__52848),
            .I(N__52845));
    Span4Mux_h I__12346 (
            .O(N__52845),
            .I(N__52842));
    Span4Mux_h I__12345 (
            .O(N__52842),
            .I(N__52839));
    Odrv4 I__12344 (
            .O(N__52839),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__12343 (
            .O(N__52836),
            .I(N__52833));
    LocalMux I__12342 (
            .O(N__52833),
            .I(N__52830));
    Odrv4 I__12341 (
            .O(N__52830),
            .I(pwm_duty_input_9));
    InMux I__12340 (
            .O(N__52827),
            .I(N__52822));
    CascadeMux I__12339 (
            .O(N__52826),
            .I(N__52819));
    InMux I__12338 (
            .O(N__52825),
            .I(N__52816));
    LocalMux I__12337 (
            .O(N__52822),
            .I(N__52813));
    InMux I__12336 (
            .O(N__52819),
            .I(N__52810));
    LocalMux I__12335 (
            .O(N__52816),
            .I(N__52807));
    Span4Mux_v I__12334 (
            .O(N__52813),
            .I(N__52804));
    LocalMux I__12333 (
            .O(N__52810),
            .I(N__52799));
    Sp12to4 I__12332 (
            .O(N__52807),
            .I(N__52799));
    Sp12to4 I__12331 (
            .O(N__52804),
            .I(N__52794));
    Span12Mux_s11_v I__12330 (
            .O(N__52799),
            .I(N__52794));
    Odrv12 I__12329 (
            .O(N__52794),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__12328 (
            .O(N__52791),
            .I(N__52788));
    LocalMux I__12327 (
            .O(N__52788),
            .I(N__52785));
    Odrv4 I__12326 (
            .O(N__52785),
            .I(pwm_duty_input_6));
    CascadeMux I__12325 (
            .O(N__52782),
            .I(N__52778));
    CascadeMux I__12324 (
            .O(N__52781),
            .I(N__52775));
    InMux I__12323 (
            .O(N__52778),
            .I(N__52771));
    InMux I__12322 (
            .O(N__52775),
            .I(N__52768));
    InMux I__12321 (
            .O(N__52774),
            .I(N__52765));
    LocalMux I__12320 (
            .O(N__52771),
            .I(N__52762));
    LocalMux I__12319 (
            .O(N__52768),
            .I(N__52757));
    LocalMux I__12318 (
            .O(N__52765),
            .I(N__52757));
    Span4Mux_v I__12317 (
            .O(N__52762),
            .I(N__52754));
    Span4Mux_v I__12316 (
            .O(N__52757),
            .I(N__52751));
    Sp12to4 I__12315 (
            .O(N__52754),
            .I(N__52746));
    Sp12to4 I__12314 (
            .O(N__52751),
            .I(N__52746));
    Odrv12 I__12313 (
            .O(N__52746),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__12312 (
            .O(N__52743),
            .I(N__52740));
    LocalMux I__12311 (
            .O(N__52740),
            .I(N__52737));
    Span4Mux_v I__12310 (
            .O(N__52737),
            .I(N__52734));
    Odrv4 I__12309 (
            .O(N__52734),
            .I(pwm_duty_input_5));
    InMux I__12308 (
            .O(N__52731),
            .I(N__52728));
    LocalMux I__12307 (
            .O(N__52728),
            .I(N__52723));
    InMux I__12306 (
            .O(N__52727),
            .I(N__52720));
    InMux I__12305 (
            .O(N__52726),
            .I(N__52717));
    Span4Mux_s3_h I__12304 (
            .O(N__52723),
            .I(N__52710));
    LocalMux I__12303 (
            .O(N__52720),
            .I(N__52710));
    LocalMux I__12302 (
            .O(N__52717),
            .I(N__52710));
    Span4Mux_v I__12301 (
            .O(N__52710),
            .I(N__52707));
    Sp12to4 I__12300 (
            .O(N__52707),
            .I(N__52704));
    Odrv12 I__12299 (
            .O(N__52704),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__12298 (
            .O(N__52701),
            .I(N__52698));
    LocalMux I__12297 (
            .O(N__52698),
            .I(N__52695));
    Odrv4 I__12296 (
            .O(N__52695),
            .I(pwm_duty_input_8));
    InMux I__12295 (
            .O(N__52692),
            .I(N__52684));
    InMux I__12294 (
            .O(N__52691),
            .I(N__52673));
    InMux I__12293 (
            .O(N__52690),
            .I(N__52673));
    InMux I__12292 (
            .O(N__52689),
            .I(N__52673));
    InMux I__12291 (
            .O(N__52688),
            .I(N__52673));
    InMux I__12290 (
            .O(N__52687),
            .I(N__52673));
    LocalMux I__12289 (
            .O(N__52684),
            .I(N__52669));
    LocalMux I__12288 (
            .O(N__52673),
            .I(N__52666));
    InMux I__12287 (
            .O(N__52672),
            .I(N__52663));
    Span4Mux_s1_h I__12286 (
            .O(N__52669),
            .I(N__52656));
    Span4Mux_v I__12285 (
            .O(N__52666),
            .I(N__52656));
    LocalMux I__12284 (
            .O(N__52663),
            .I(N__52656));
    Span4Mux_h I__12283 (
            .O(N__52656),
            .I(N__52653));
    Odrv4 I__12282 (
            .O(N__52653),
            .I(\current_shift_inst.PI_CTRL.N_150 ));
    InMux I__12281 (
            .O(N__52650),
            .I(N__52635));
    InMux I__12280 (
            .O(N__52649),
            .I(N__52635));
    InMux I__12279 (
            .O(N__52648),
            .I(N__52635));
    InMux I__12278 (
            .O(N__52647),
            .I(N__52635));
    InMux I__12277 (
            .O(N__52646),
            .I(N__52635));
    LocalMux I__12276 (
            .O(N__52635),
            .I(N__52631));
    InMux I__12275 (
            .O(N__52634),
            .I(N__52628));
    Span4Mux_v I__12274 (
            .O(N__52631),
            .I(N__52621));
    LocalMux I__12273 (
            .O(N__52628),
            .I(N__52618));
    InMux I__12272 (
            .O(N__52627),
            .I(N__52609));
    InMux I__12271 (
            .O(N__52626),
            .I(N__52609));
    InMux I__12270 (
            .O(N__52625),
            .I(N__52609));
    InMux I__12269 (
            .O(N__52624),
            .I(N__52609));
    Span4Mux_h I__12268 (
            .O(N__52621),
            .I(N__52606));
    Span4Mux_v I__12267 (
            .O(N__52618),
            .I(N__52603));
    LocalMux I__12266 (
            .O(N__52609),
            .I(N__52600));
    Sp12to4 I__12265 (
            .O(N__52606),
            .I(N__52593));
    Sp12to4 I__12264 (
            .O(N__52603),
            .I(N__52593));
    Span12Mux_s4_h I__12263 (
            .O(N__52600),
            .I(N__52593));
    Odrv12 I__12262 (
            .O(N__52593),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__12261 (
            .O(N__52590),
            .I(N__52583));
    CascadeMux I__12260 (
            .O(N__52589),
            .I(N__52580));
    CascadeMux I__12259 (
            .O(N__52588),
            .I(N__52577));
    InMux I__12258 (
            .O(N__52587),
            .I(N__52566));
    InMux I__12257 (
            .O(N__52586),
            .I(N__52566));
    InMux I__12256 (
            .O(N__52583),
            .I(N__52566));
    InMux I__12255 (
            .O(N__52580),
            .I(N__52566));
    InMux I__12254 (
            .O(N__52577),
            .I(N__52566));
    LocalMux I__12253 (
            .O(N__52566),
            .I(N__52563));
    Span4Mux_v I__12252 (
            .O(N__52563),
            .I(N__52557));
    InMux I__12251 (
            .O(N__52562),
            .I(N__52552));
    InMux I__12250 (
            .O(N__52561),
            .I(N__52552));
    InMux I__12249 (
            .O(N__52560),
            .I(N__52549));
    Sp12to4 I__12248 (
            .O(N__52557),
            .I(N__52542));
    LocalMux I__12247 (
            .O(N__52552),
            .I(N__52542));
    LocalMux I__12246 (
            .O(N__52549),
            .I(N__52542));
    Span12Mux_s9_h I__12245 (
            .O(N__52542),
            .I(N__52539));
    Odrv12 I__12244 (
            .O(N__52539),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_11 ));
    InMux I__12243 (
            .O(N__52536),
            .I(N__52533));
    LocalMux I__12242 (
            .O(N__52533),
            .I(N__52528));
    InMux I__12241 (
            .O(N__52532),
            .I(N__52523));
    InMux I__12240 (
            .O(N__52531),
            .I(N__52523));
    Span4Mux_s3_h I__12239 (
            .O(N__52528),
            .I(N__52518));
    LocalMux I__12238 (
            .O(N__52523),
            .I(N__52518));
    Span4Mux_v I__12237 (
            .O(N__52518),
            .I(N__52515));
    Sp12to4 I__12236 (
            .O(N__52515),
            .I(N__52512));
    Odrv12 I__12235 (
            .O(N__52512),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__12234 (
            .O(N__52509),
            .I(N__52506));
    LocalMux I__12233 (
            .O(N__52506),
            .I(N__52503));
    Odrv4 I__12232 (
            .O(N__52503),
            .I(pwm_duty_input_7));
    ClkMux I__12231 (
            .O(N__52500),
            .I(N__52092));
    ClkMux I__12230 (
            .O(N__52499),
            .I(N__52092));
    ClkMux I__12229 (
            .O(N__52498),
            .I(N__52092));
    ClkMux I__12228 (
            .O(N__52497),
            .I(N__52092));
    ClkMux I__12227 (
            .O(N__52496),
            .I(N__52092));
    ClkMux I__12226 (
            .O(N__52495),
            .I(N__52092));
    ClkMux I__12225 (
            .O(N__52494),
            .I(N__52092));
    ClkMux I__12224 (
            .O(N__52493),
            .I(N__52092));
    ClkMux I__12223 (
            .O(N__52492),
            .I(N__52092));
    ClkMux I__12222 (
            .O(N__52491),
            .I(N__52092));
    ClkMux I__12221 (
            .O(N__52490),
            .I(N__52092));
    ClkMux I__12220 (
            .O(N__52489),
            .I(N__52092));
    ClkMux I__12219 (
            .O(N__52488),
            .I(N__52092));
    ClkMux I__12218 (
            .O(N__52487),
            .I(N__52092));
    ClkMux I__12217 (
            .O(N__52486),
            .I(N__52092));
    ClkMux I__12216 (
            .O(N__52485),
            .I(N__52092));
    ClkMux I__12215 (
            .O(N__52484),
            .I(N__52092));
    ClkMux I__12214 (
            .O(N__52483),
            .I(N__52092));
    ClkMux I__12213 (
            .O(N__52482),
            .I(N__52092));
    ClkMux I__12212 (
            .O(N__52481),
            .I(N__52092));
    ClkMux I__12211 (
            .O(N__52480),
            .I(N__52092));
    ClkMux I__12210 (
            .O(N__52479),
            .I(N__52092));
    ClkMux I__12209 (
            .O(N__52478),
            .I(N__52092));
    ClkMux I__12208 (
            .O(N__52477),
            .I(N__52092));
    ClkMux I__12207 (
            .O(N__52476),
            .I(N__52092));
    ClkMux I__12206 (
            .O(N__52475),
            .I(N__52092));
    ClkMux I__12205 (
            .O(N__52474),
            .I(N__52092));
    ClkMux I__12204 (
            .O(N__52473),
            .I(N__52092));
    ClkMux I__12203 (
            .O(N__52472),
            .I(N__52092));
    ClkMux I__12202 (
            .O(N__52471),
            .I(N__52092));
    ClkMux I__12201 (
            .O(N__52470),
            .I(N__52092));
    ClkMux I__12200 (
            .O(N__52469),
            .I(N__52092));
    ClkMux I__12199 (
            .O(N__52468),
            .I(N__52092));
    ClkMux I__12198 (
            .O(N__52467),
            .I(N__52092));
    ClkMux I__12197 (
            .O(N__52466),
            .I(N__52092));
    ClkMux I__12196 (
            .O(N__52465),
            .I(N__52092));
    ClkMux I__12195 (
            .O(N__52464),
            .I(N__52092));
    ClkMux I__12194 (
            .O(N__52463),
            .I(N__52092));
    ClkMux I__12193 (
            .O(N__52462),
            .I(N__52092));
    ClkMux I__12192 (
            .O(N__52461),
            .I(N__52092));
    ClkMux I__12191 (
            .O(N__52460),
            .I(N__52092));
    ClkMux I__12190 (
            .O(N__52459),
            .I(N__52092));
    ClkMux I__12189 (
            .O(N__52458),
            .I(N__52092));
    ClkMux I__12188 (
            .O(N__52457),
            .I(N__52092));
    ClkMux I__12187 (
            .O(N__52456),
            .I(N__52092));
    ClkMux I__12186 (
            .O(N__52455),
            .I(N__52092));
    ClkMux I__12185 (
            .O(N__52454),
            .I(N__52092));
    ClkMux I__12184 (
            .O(N__52453),
            .I(N__52092));
    ClkMux I__12183 (
            .O(N__52452),
            .I(N__52092));
    ClkMux I__12182 (
            .O(N__52451),
            .I(N__52092));
    ClkMux I__12181 (
            .O(N__52450),
            .I(N__52092));
    ClkMux I__12180 (
            .O(N__52449),
            .I(N__52092));
    ClkMux I__12179 (
            .O(N__52448),
            .I(N__52092));
    ClkMux I__12178 (
            .O(N__52447),
            .I(N__52092));
    ClkMux I__12177 (
            .O(N__52446),
            .I(N__52092));
    ClkMux I__12176 (
            .O(N__52445),
            .I(N__52092));
    ClkMux I__12175 (
            .O(N__52444),
            .I(N__52092));
    ClkMux I__12174 (
            .O(N__52443),
            .I(N__52092));
    ClkMux I__12173 (
            .O(N__52442),
            .I(N__52092));
    ClkMux I__12172 (
            .O(N__52441),
            .I(N__52092));
    ClkMux I__12171 (
            .O(N__52440),
            .I(N__52092));
    ClkMux I__12170 (
            .O(N__52439),
            .I(N__52092));
    ClkMux I__12169 (
            .O(N__52438),
            .I(N__52092));
    ClkMux I__12168 (
            .O(N__52437),
            .I(N__52092));
    ClkMux I__12167 (
            .O(N__52436),
            .I(N__52092));
    ClkMux I__12166 (
            .O(N__52435),
            .I(N__52092));
    ClkMux I__12165 (
            .O(N__52434),
            .I(N__52092));
    ClkMux I__12164 (
            .O(N__52433),
            .I(N__52092));
    ClkMux I__12163 (
            .O(N__52432),
            .I(N__52092));
    ClkMux I__12162 (
            .O(N__52431),
            .I(N__52092));
    ClkMux I__12161 (
            .O(N__52430),
            .I(N__52092));
    ClkMux I__12160 (
            .O(N__52429),
            .I(N__52092));
    ClkMux I__12159 (
            .O(N__52428),
            .I(N__52092));
    ClkMux I__12158 (
            .O(N__52427),
            .I(N__52092));
    ClkMux I__12157 (
            .O(N__52426),
            .I(N__52092));
    ClkMux I__12156 (
            .O(N__52425),
            .I(N__52092));
    ClkMux I__12155 (
            .O(N__52424),
            .I(N__52092));
    ClkMux I__12154 (
            .O(N__52423),
            .I(N__52092));
    ClkMux I__12153 (
            .O(N__52422),
            .I(N__52092));
    ClkMux I__12152 (
            .O(N__52421),
            .I(N__52092));
    ClkMux I__12151 (
            .O(N__52420),
            .I(N__52092));
    ClkMux I__12150 (
            .O(N__52419),
            .I(N__52092));
    ClkMux I__12149 (
            .O(N__52418),
            .I(N__52092));
    ClkMux I__12148 (
            .O(N__52417),
            .I(N__52092));
    ClkMux I__12147 (
            .O(N__52416),
            .I(N__52092));
    ClkMux I__12146 (
            .O(N__52415),
            .I(N__52092));
    ClkMux I__12145 (
            .O(N__52414),
            .I(N__52092));
    ClkMux I__12144 (
            .O(N__52413),
            .I(N__52092));
    ClkMux I__12143 (
            .O(N__52412),
            .I(N__52092));
    ClkMux I__12142 (
            .O(N__52411),
            .I(N__52092));
    ClkMux I__12141 (
            .O(N__52410),
            .I(N__52092));
    ClkMux I__12140 (
            .O(N__52409),
            .I(N__52092));
    ClkMux I__12139 (
            .O(N__52408),
            .I(N__52092));
    ClkMux I__12138 (
            .O(N__52407),
            .I(N__52092));
    ClkMux I__12137 (
            .O(N__52406),
            .I(N__52092));
    ClkMux I__12136 (
            .O(N__52405),
            .I(N__52092));
    ClkMux I__12135 (
            .O(N__52404),
            .I(N__52092));
    ClkMux I__12134 (
            .O(N__52403),
            .I(N__52092));
    ClkMux I__12133 (
            .O(N__52402),
            .I(N__52092));
    ClkMux I__12132 (
            .O(N__52401),
            .I(N__52092));
    ClkMux I__12131 (
            .O(N__52400),
            .I(N__52092));
    ClkMux I__12130 (
            .O(N__52399),
            .I(N__52092));
    ClkMux I__12129 (
            .O(N__52398),
            .I(N__52092));
    ClkMux I__12128 (
            .O(N__52397),
            .I(N__52092));
    ClkMux I__12127 (
            .O(N__52396),
            .I(N__52092));
    ClkMux I__12126 (
            .O(N__52395),
            .I(N__52092));
    ClkMux I__12125 (
            .O(N__52394),
            .I(N__52092));
    ClkMux I__12124 (
            .O(N__52393),
            .I(N__52092));
    ClkMux I__12123 (
            .O(N__52392),
            .I(N__52092));
    ClkMux I__12122 (
            .O(N__52391),
            .I(N__52092));
    ClkMux I__12121 (
            .O(N__52390),
            .I(N__52092));
    ClkMux I__12120 (
            .O(N__52389),
            .I(N__52092));
    ClkMux I__12119 (
            .O(N__52388),
            .I(N__52092));
    ClkMux I__12118 (
            .O(N__52387),
            .I(N__52092));
    ClkMux I__12117 (
            .O(N__52386),
            .I(N__52092));
    ClkMux I__12116 (
            .O(N__52385),
            .I(N__52092));
    ClkMux I__12115 (
            .O(N__52384),
            .I(N__52092));
    ClkMux I__12114 (
            .O(N__52383),
            .I(N__52092));
    ClkMux I__12113 (
            .O(N__52382),
            .I(N__52092));
    ClkMux I__12112 (
            .O(N__52381),
            .I(N__52092));
    ClkMux I__12111 (
            .O(N__52380),
            .I(N__52092));
    ClkMux I__12110 (
            .O(N__52379),
            .I(N__52092));
    ClkMux I__12109 (
            .O(N__52378),
            .I(N__52092));
    ClkMux I__12108 (
            .O(N__52377),
            .I(N__52092));
    ClkMux I__12107 (
            .O(N__52376),
            .I(N__52092));
    ClkMux I__12106 (
            .O(N__52375),
            .I(N__52092));
    ClkMux I__12105 (
            .O(N__52374),
            .I(N__52092));
    ClkMux I__12104 (
            .O(N__52373),
            .I(N__52092));
    ClkMux I__12103 (
            .O(N__52372),
            .I(N__52092));
    ClkMux I__12102 (
            .O(N__52371),
            .I(N__52092));
    ClkMux I__12101 (
            .O(N__52370),
            .I(N__52092));
    ClkMux I__12100 (
            .O(N__52369),
            .I(N__52092));
    ClkMux I__12099 (
            .O(N__52368),
            .I(N__52092));
    ClkMux I__12098 (
            .O(N__52367),
            .I(N__52092));
    ClkMux I__12097 (
            .O(N__52366),
            .I(N__52092));
    ClkMux I__12096 (
            .O(N__52365),
            .I(N__52092));
    GlobalMux I__12095 (
            .O(N__52092),
            .I(clk_100mhz_0));
    InMux I__12094 (
            .O(N__52089),
            .I(N__52079));
    InMux I__12093 (
            .O(N__52088),
            .I(N__52076));
    InMux I__12092 (
            .O(N__52087),
            .I(N__52073));
    InMux I__12091 (
            .O(N__52086),
            .I(N__52070));
    InMux I__12090 (
            .O(N__52085),
            .I(N__52067));
    InMux I__12089 (
            .O(N__52084),
            .I(N__52064));
    InMux I__12088 (
            .O(N__52083),
            .I(N__52061));
    InMux I__12087 (
            .O(N__52082),
            .I(N__52058));
    LocalMux I__12086 (
            .O(N__52079),
            .I(N__52055));
    LocalMux I__12085 (
            .O(N__52076),
            .I(N__52052));
    LocalMux I__12084 (
            .O(N__52073),
            .I(N__52049));
    LocalMux I__12083 (
            .O(N__52070),
            .I(N__52027));
    LocalMux I__12082 (
            .O(N__52067),
            .I(N__51983));
    LocalMux I__12081 (
            .O(N__52064),
            .I(N__51948));
    LocalMux I__12080 (
            .O(N__52061),
            .I(N__51936));
    LocalMux I__12079 (
            .O(N__52058),
            .I(N__51929));
    Glb2LocalMux I__12078 (
            .O(N__52055),
            .I(N__51699));
    Glb2LocalMux I__12077 (
            .O(N__52052),
            .I(N__51699));
    Glb2LocalMux I__12076 (
            .O(N__52049),
            .I(N__51699));
    SRMux I__12075 (
            .O(N__52048),
            .I(N__51699));
    SRMux I__12074 (
            .O(N__52047),
            .I(N__51699));
    SRMux I__12073 (
            .O(N__52046),
            .I(N__51699));
    SRMux I__12072 (
            .O(N__52045),
            .I(N__51699));
    SRMux I__12071 (
            .O(N__52044),
            .I(N__51699));
    SRMux I__12070 (
            .O(N__52043),
            .I(N__51699));
    SRMux I__12069 (
            .O(N__52042),
            .I(N__51699));
    SRMux I__12068 (
            .O(N__52041),
            .I(N__51699));
    SRMux I__12067 (
            .O(N__52040),
            .I(N__51699));
    SRMux I__12066 (
            .O(N__52039),
            .I(N__51699));
    SRMux I__12065 (
            .O(N__52038),
            .I(N__51699));
    SRMux I__12064 (
            .O(N__52037),
            .I(N__51699));
    SRMux I__12063 (
            .O(N__52036),
            .I(N__51699));
    SRMux I__12062 (
            .O(N__52035),
            .I(N__51699));
    SRMux I__12061 (
            .O(N__52034),
            .I(N__51699));
    SRMux I__12060 (
            .O(N__52033),
            .I(N__51699));
    SRMux I__12059 (
            .O(N__52032),
            .I(N__51699));
    SRMux I__12058 (
            .O(N__52031),
            .I(N__51699));
    SRMux I__12057 (
            .O(N__52030),
            .I(N__51699));
    Glb2LocalMux I__12056 (
            .O(N__52027),
            .I(N__51699));
    SRMux I__12055 (
            .O(N__52026),
            .I(N__51699));
    SRMux I__12054 (
            .O(N__52025),
            .I(N__51699));
    SRMux I__12053 (
            .O(N__52024),
            .I(N__51699));
    SRMux I__12052 (
            .O(N__52023),
            .I(N__51699));
    SRMux I__12051 (
            .O(N__52022),
            .I(N__51699));
    SRMux I__12050 (
            .O(N__52021),
            .I(N__51699));
    SRMux I__12049 (
            .O(N__52020),
            .I(N__51699));
    SRMux I__12048 (
            .O(N__52019),
            .I(N__51699));
    SRMux I__12047 (
            .O(N__52018),
            .I(N__51699));
    SRMux I__12046 (
            .O(N__52017),
            .I(N__51699));
    SRMux I__12045 (
            .O(N__52016),
            .I(N__51699));
    SRMux I__12044 (
            .O(N__52015),
            .I(N__51699));
    SRMux I__12043 (
            .O(N__52014),
            .I(N__51699));
    SRMux I__12042 (
            .O(N__52013),
            .I(N__51699));
    SRMux I__12041 (
            .O(N__52012),
            .I(N__51699));
    SRMux I__12040 (
            .O(N__52011),
            .I(N__51699));
    SRMux I__12039 (
            .O(N__52010),
            .I(N__51699));
    SRMux I__12038 (
            .O(N__52009),
            .I(N__51699));
    SRMux I__12037 (
            .O(N__52008),
            .I(N__51699));
    SRMux I__12036 (
            .O(N__52007),
            .I(N__51699));
    SRMux I__12035 (
            .O(N__52006),
            .I(N__51699));
    SRMux I__12034 (
            .O(N__52005),
            .I(N__51699));
    SRMux I__12033 (
            .O(N__52004),
            .I(N__51699));
    SRMux I__12032 (
            .O(N__52003),
            .I(N__51699));
    SRMux I__12031 (
            .O(N__52002),
            .I(N__51699));
    SRMux I__12030 (
            .O(N__52001),
            .I(N__51699));
    SRMux I__12029 (
            .O(N__52000),
            .I(N__51699));
    SRMux I__12028 (
            .O(N__51999),
            .I(N__51699));
    SRMux I__12027 (
            .O(N__51998),
            .I(N__51699));
    SRMux I__12026 (
            .O(N__51997),
            .I(N__51699));
    SRMux I__12025 (
            .O(N__51996),
            .I(N__51699));
    SRMux I__12024 (
            .O(N__51995),
            .I(N__51699));
    SRMux I__12023 (
            .O(N__51994),
            .I(N__51699));
    SRMux I__12022 (
            .O(N__51993),
            .I(N__51699));
    SRMux I__12021 (
            .O(N__51992),
            .I(N__51699));
    SRMux I__12020 (
            .O(N__51991),
            .I(N__51699));
    SRMux I__12019 (
            .O(N__51990),
            .I(N__51699));
    SRMux I__12018 (
            .O(N__51989),
            .I(N__51699));
    SRMux I__12017 (
            .O(N__51988),
            .I(N__51699));
    SRMux I__12016 (
            .O(N__51987),
            .I(N__51699));
    SRMux I__12015 (
            .O(N__51986),
            .I(N__51699));
    Glb2LocalMux I__12014 (
            .O(N__51983),
            .I(N__51699));
    SRMux I__12013 (
            .O(N__51982),
            .I(N__51699));
    SRMux I__12012 (
            .O(N__51981),
            .I(N__51699));
    SRMux I__12011 (
            .O(N__51980),
            .I(N__51699));
    SRMux I__12010 (
            .O(N__51979),
            .I(N__51699));
    SRMux I__12009 (
            .O(N__51978),
            .I(N__51699));
    SRMux I__12008 (
            .O(N__51977),
            .I(N__51699));
    SRMux I__12007 (
            .O(N__51976),
            .I(N__51699));
    SRMux I__12006 (
            .O(N__51975),
            .I(N__51699));
    SRMux I__12005 (
            .O(N__51974),
            .I(N__51699));
    SRMux I__12004 (
            .O(N__51973),
            .I(N__51699));
    SRMux I__12003 (
            .O(N__51972),
            .I(N__51699));
    SRMux I__12002 (
            .O(N__51971),
            .I(N__51699));
    SRMux I__12001 (
            .O(N__51970),
            .I(N__51699));
    SRMux I__12000 (
            .O(N__51969),
            .I(N__51699));
    SRMux I__11999 (
            .O(N__51968),
            .I(N__51699));
    SRMux I__11998 (
            .O(N__51967),
            .I(N__51699));
    SRMux I__11997 (
            .O(N__51966),
            .I(N__51699));
    SRMux I__11996 (
            .O(N__51965),
            .I(N__51699));
    SRMux I__11995 (
            .O(N__51964),
            .I(N__51699));
    SRMux I__11994 (
            .O(N__51963),
            .I(N__51699));
    SRMux I__11993 (
            .O(N__51962),
            .I(N__51699));
    SRMux I__11992 (
            .O(N__51961),
            .I(N__51699));
    SRMux I__11991 (
            .O(N__51960),
            .I(N__51699));
    SRMux I__11990 (
            .O(N__51959),
            .I(N__51699));
    SRMux I__11989 (
            .O(N__51958),
            .I(N__51699));
    SRMux I__11988 (
            .O(N__51957),
            .I(N__51699));
    SRMux I__11987 (
            .O(N__51956),
            .I(N__51699));
    SRMux I__11986 (
            .O(N__51955),
            .I(N__51699));
    SRMux I__11985 (
            .O(N__51954),
            .I(N__51699));
    SRMux I__11984 (
            .O(N__51953),
            .I(N__51699));
    SRMux I__11983 (
            .O(N__51952),
            .I(N__51699));
    SRMux I__11982 (
            .O(N__51951),
            .I(N__51699));
    Glb2LocalMux I__11981 (
            .O(N__51948),
            .I(N__51699));
    SRMux I__11980 (
            .O(N__51947),
            .I(N__51699));
    SRMux I__11979 (
            .O(N__51946),
            .I(N__51699));
    SRMux I__11978 (
            .O(N__51945),
            .I(N__51699));
    SRMux I__11977 (
            .O(N__51944),
            .I(N__51699));
    SRMux I__11976 (
            .O(N__51943),
            .I(N__51699));
    SRMux I__11975 (
            .O(N__51942),
            .I(N__51699));
    SRMux I__11974 (
            .O(N__51941),
            .I(N__51699));
    SRMux I__11973 (
            .O(N__51940),
            .I(N__51699));
    SRMux I__11972 (
            .O(N__51939),
            .I(N__51699));
    Glb2LocalMux I__11971 (
            .O(N__51936),
            .I(N__51699));
    SRMux I__11970 (
            .O(N__51935),
            .I(N__51699));
    SRMux I__11969 (
            .O(N__51934),
            .I(N__51699));
    SRMux I__11968 (
            .O(N__51933),
            .I(N__51699));
    SRMux I__11967 (
            .O(N__51932),
            .I(N__51699));
    Glb2LocalMux I__11966 (
            .O(N__51929),
            .I(N__51699));
    SRMux I__11965 (
            .O(N__51928),
            .I(N__51699));
    GlobalMux I__11964 (
            .O(N__51699),
            .I(N__51696));
    gio2CtrlBuf I__11963 (
            .O(N__51696),
            .I(red_c_g));
    InMux I__11962 (
            .O(N__51693),
            .I(N__51690));
    LocalMux I__11961 (
            .O(N__51690),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    CascadeMux I__11960 (
            .O(N__51687),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    InMux I__11959 (
            .O(N__51684),
            .I(N__51681));
    LocalMux I__11958 (
            .O(N__51681),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__11957 (
            .O(N__51678),
            .I(N__51669));
    InMux I__11956 (
            .O(N__51677),
            .I(N__51669));
    InMux I__11955 (
            .O(N__51676),
            .I(N__51669));
    LocalMux I__11954 (
            .O(N__51669),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__11953 (
            .O(N__51666),
            .I(N__51663));
    LocalMux I__11952 (
            .O(N__51663),
            .I(N__51660));
    Span12Mux_v I__11951 (
            .O(N__51660),
            .I(N__51657));
    Span12Mux_h I__11950 (
            .O(N__51657),
            .I(N__51654));
    Odrv12 I__11949 (
            .O(N__51654),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__11948 (
            .O(N__51651),
            .I(N__51648));
    LocalMux I__11947 (
            .O(N__51648),
            .I(N__51645));
    Span4Mux_v I__11946 (
            .O(N__51645),
            .I(N__51642));
    Span4Mux_h I__11945 (
            .O(N__51642),
            .I(N__51639));
    Sp12to4 I__11944 (
            .O(N__51639),
            .I(N__51636));
    Odrv12 I__11943 (
            .O(N__51636),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__11942 (
            .O(N__51633),
            .I(N__51630));
    LocalMux I__11941 (
            .O(N__51630),
            .I(N__51627));
    Span4Mux_v I__11940 (
            .O(N__51627),
            .I(N__51624));
    Odrv4 I__11939 (
            .O(N__51624),
            .I(pwm_duty_input_2));
    InMux I__11938 (
            .O(N__51621),
            .I(N__51618));
    LocalMux I__11937 (
            .O(N__51618),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__11936 (
            .O(N__51615),
            .I(N__51612));
    LocalMux I__11935 (
            .O(N__51612),
            .I(N__51609));
    Odrv4 I__11934 (
            .O(N__51609),
            .I(pwm_duty_input_0));
    InMux I__11933 (
            .O(N__51606),
            .I(N__51597));
    InMux I__11932 (
            .O(N__51605),
            .I(N__51597));
    InMux I__11931 (
            .O(N__51604),
            .I(N__51597));
    LocalMux I__11930 (
            .O(N__51597),
            .I(\current_shift_inst.PI_CTRL.N_152 ));
    InMux I__11929 (
            .O(N__51594),
            .I(N__51591));
    LocalMux I__11928 (
            .O(N__51591),
            .I(N__51588));
    Span4Mux_v I__11927 (
            .O(N__51588),
            .I(N__51585));
    Sp12to4 I__11926 (
            .O(N__51585),
            .I(N__51582));
    Span12Mux_h I__11925 (
            .O(N__51582),
            .I(N__51579));
    Odrv12 I__11924 (
            .O(N__51579),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__11923 (
            .O(N__51576),
            .I(N__51573));
    LocalMux I__11922 (
            .O(N__51573),
            .I(N__51570));
    Odrv4 I__11921 (
            .O(N__51570),
            .I(pwm_duty_input_1));
    InMux I__11920 (
            .O(N__51567),
            .I(N__51564));
    LocalMux I__11919 (
            .O(N__51564),
            .I(N__51559));
    InMux I__11918 (
            .O(N__51563),
            .I(N__51556));
    InMux I__11917 (
            .O(N__51562),
            .I(N__51553));
    Span4Mux_v I__11916 (
            .O(N__51559),
            .I(N__51550));
    LocalMux I__11915 (
            .O(N__51556),
            .I(N__51545));
    LocalMux I__11914 (
            .O(N__51553),
            .I(N__51545));
    Sp12to4 I__11913 (
            .O(N__51550),
            .I(N__51542));
    Span12Mux_v I__11912 (
            .O(N__51545),
            .I(N__51539));
    Span12Mux_s8_h I__11911 (
            .O(N__51542),
            .I(N__51536));
    Span12Mux_h I__11910 (
            .O(N__51539),
            .I(N__51533));
    Odrv12 I__11909 (
            .O(N__51536),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv12 I__11908 (
            .O(N__51533),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__11907 (
            .O(N__51528),
            .I(N__51524));
    InMux I__11906 (
            .O(N__51527),
            .I(N__51521));
    LocalMux I__11905 (
            .O(N__51524),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__11904 (
            .O(N__51521),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__11903 (
            .O(N__51516),
            .I(N__51513));
    LocalMux I__11902 (
            .O(N__51513),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__11901 (
            .O(N__51510),
            .I(N__51507));
    LocalMux I__11900 (
            .O(N__51507),
            .I(N__51504));
    Span4Mux_s0_h I__11899 (
            .O(N__51504),
            .I(N__51501));
    Odrv4 I__11898 (
            .O(N__51501),
            .I(pwm_duty_input_3));
    CascadeMux I__11897 (
            .O(N__51498),
            .I(N__51493));
    InMux I__11896 (
            .O(N__51497),
            .I(N__51490));
    InMux I__11895 (
            .O(N__51496),
            .I(N__51487));
    InMux I__11894 (
            .O(N__51493),
            .I(N__51484));
    LocalMux I__11893 (
            .O(N__51490),
            .I(N__51481));
    LocalMux I__11892 (
            .O(N__51487),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__11891 (
            .O(N__51484),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv12 I__11890 (
            .O(N__51481),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__11889 (
            .O(N__51474),
            .I(N__51471));
    LocalMux I__11888 (
            .O(N__51471),
            .I(N__51468));
    Odrv4 I__11887 (
            .O(N__51468),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__11886 (
            .O(N__51465),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__11885 (
            .O(N__51462),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__11884 (
            .O(N__51459),
            .I(N__51456));
    LocalMux I__11883 (
            .O(N__51456),
            .I(N__51453));
    Odrv4 I__11882 (
            .O(N__51453),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__11881 (
            .O(N__51450),
            .I(N__51446));
    InMux I__11880 (
            .O(N__51449),
            .I(N__51443));
    LocalMux I__11879 (
            .O(N__51446),
            .I(N__51440));
    LocalMux I__11878 (
            .O(N__51443),
            .I(N__51437));
    Span12Mux_h I__11877 (
            .O(N__51440),
            .I(N__51434));
    Span4Mux_v I__11876 (
            .O(N__51437),
            .I(N__51431));
    Odrv12 I__11875 (
            .O(N__51434),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__11874 (
            .O(N__51431),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__11873 (
            .O(N__51426),
            .I(N__51422));
    InMux I__11872 (
            .O(N__51425),
            .I(N__51418));
    LocalMux I__11871 (
            .O(N__51422),
            .I(N__51415));
    InMux I__11870 (
            .O(N__51421),
            .I(N__51412));
    LocalMux I__11869 (
            .O(N__51418),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv12 I__11868 (
            .O(N__51415),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    LocalMux I__11867 (
            .O(N__51412),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__11866 (
            .O(N__51405),
            .I(N__51402));
    LocalMux I__11865 (
            .O(N__51402),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ));
    InMux I__11864 (
            .O(N__51399),
            .I(N__51396));
    LocalMux I__11863 (
            .O(N__51396),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ));
    InMux I__11862 (
            .O(N__51393),
            .I(N__51390));
    LocalMux I__11861 (
            .O(N__51390),
            .I(N__51387));
    Odrv12 I__11860 (
            .O(N__51387),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__11859 (
            .O(N__51384),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    CascadeMux I__11858 (
            .O(N__51381),
            .I(N__51375));
    InMux I__11857 (
            .O(N__51380),
            .I(N__51371));
    CascadeMux I__11856 (
            .O(N__51379),
            .I(N__51364));
    CascadeMux I__11855 (
            .O(N__51378),
            .I(N__51361));
    InMux I__11854 (
            .O(N__51375),
            .I(N__51355));
    InMux I__11853 (
            .O(N__51374),
            .I(N__51352));
    LocalMux I__11852 (
            .O(N__51371),
            .I(N__51349));
    InMux I__11851 (
            .O(N__51370),
            .I(N__51346));
    InMux I__11850 (
            .O(N__51369),
            .I(N__51337));
    InMux I__11849 (
            .O(N__51368),
            .I(N__51337));
    InMux I__11848 (
            .O(N__51367),
            .I(N__51337));
    InMux I__11847 (
            .O(N__51364),
            .I(N__51337));
    InMux I__11846 (
            .O(N__51361),
            .I(N__51328));
    InMux I__11845 (
            .O(N__51360),
            .I(N__51328));
    InMux I__11844 (
            .O(N__51359),
            .I(N__51328));
    InMux I__11843 (
            .O(N__51358),
            .I(N__51328));
    LocalMux I__11842 (
            .O(N__51355),
            .I(N__51323));
    LocalMux I__11841 (
            .O(N__51352),
            .I(N__51323));
    Span4Mux_h I__11840 (
            .O(N__51349),
            .I(N__51320));
    LocalMux I__11839 (
            .O(N__51346),
            .I(N__51317));
    LocalMux I__11838 (
            .O(N__51337),
            .I(N__51314));
    LocalMux I__11837 (
            .O(N__51328),
            .I(N__51309));
    Span4Mux_h I__11836 (
            .O(N__51323),
            .I(N__51309));
    Odrv4 I__11835 (
            .O(N__51320),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv12 I__11834 (
            .O(N__51317),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv12 I__11833 (
            .O(N__51314),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__11832 (
            .O(N__51309),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__11831 (
            .O(N__51300),
            .I(N__51296));
    InMux I__11830 (
            .O(N__51299),
            .I(N__51293));
    LocalMux I__11829 (
            .O(N__51296),
            .I(N__51290));
    LocalMux I__11828 (
            .O(N__51293),
            .I(N__51287));
    Span4Mux_v I__11827 (
            .O(N__51290),
            .I(N__51284));
    Span4Mux_v I__11826 (
            .O(N__51287),
            .I(N__51279));
    Span4Mux_h I__11825 (
            .O(N__51284),
            .I(N__51279));
    Span4Mux_h I__11824 (
            .O(N__51279),
            .I(N__51276));
    Odrv4 I__11823 (
            .O(N__51276),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__11822 (
            .O(N__51273),
            .I(N__51270));
    LocalMux I__11821 (
            .O(N__51270),
            .I(N__51267));
    Odrv4 I__11820 (
            .O(N__51267),
            .I(\pwm_generator_inst.un19_threshold_0_axb_1 ));
    InMux I__11819 (
            .O(N__51264),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__11818 (
            .O(N__51261),
            .I(N__51257));
    InMux I__11817 (
            .O(N__51260),
            .I(N__51254));
    LocalMux I__11816 (
            .O(N__51257),
            .I(N__51250));
    LocalMux I__11815 (
            .O(N__51254),
            .I(N__51247));
    InMux I__11814 (
            .O(N__51253),
            .I(N__51244));
    Span4Mux_v I__11813 (
            .O(N__51250),
            .I(N__51239));
    Span4Mux_h I__11812 (
            .O(N__51247),
            .I(N__51239));
    LocalMux I__11811 (
            .O(N__51244),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__11810 (
            .O(N__51239),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__11809 (
            .O(N__51234),
            .I(N__51231));
    LocalMux I__11808 (
            .O(N__51231),
            .I(N__51228));
    Odrv12 I__11807 (
            .O(N__51228),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__11806 (
            .O(N__51225),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__11805 (
            .O(N__51222),
            .I(N__51218));
    InMux I__11804 (
            .O(N__51221),
            .I(N__51215));
    LocalMux I__11803 (
            .O(N__51218),
            .I(N__51212));
    LocalMux I__11802 (
            .O(N__51215),
            .I(N__51207));
    Span4Mux_h I__11801 (
            .O(N__51212),
            .I(N__51207));
    Odrv4 I__11800 (
            .O(N__51207),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__11799 (
            .O(N__51204),
            .I(N__51201));
    LocalMux I__11798 (
            .O(N__51201),
            .I(N__51198));
    Odrv12 I__11797 (
            .O(N__51198),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__11796 (
            .O(N__51195),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__11795 (
            .O(N__51192),
            .I(N__51187));
    InMux I__11794 (
            .O(N__51191),
            .I(N__51184));
    InMux I__11793 (
            .O(N__51190),
            .I(N__51181));
    LocalMux I__11792 (
            .O(N__51187),
            .I(N__51178));
    LocalMux I__11791 (
            .O(N__51184),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__11790 (
            .O(N__51181),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv12 I__11789 (
            .O(N__51178),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__11788 (
            .O(N__51171),
            .I(N__51168));
    LocalMux I__11787 (
            .O(N__51168),
            .I(N__51165));
    Span4Mux_h I__11786 (
            .O(N__51165),
            .I(N__51162));
    Odrv4 I__11785 (
            .O(N__51162),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__11784 (
            .O(N__51159),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__11783 (
            .O(N__51156),
            .I(N__51153));
    LocalMux I__11782 (
            .O(N__51153),
            .I(N__51150));
    Span4Mux_h I__11781 (
            .O(N__51150),
            .I(N__51145));
    InMux I__11780 (
            .O(N__51149),
            .I(N__51142));
    InMux I__11779 (
            .O(N__51148),
            .I(N__51139));
    Span4Mux_h I__11778 (
            .O(N__51145),
            .I(N__51136));
    LocalMux I__11777 (
            .O(N__51142),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__11776 (
            .O(N__51139),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__11775 (
            .O(N__51136),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__11774 (
            .O(N__51129),
            .I(N__51126));
    LocalMux I__11773 (
            .O(N__51126),
            .I(N__51123));
    Odrv12 I__11772 (
            .O(N__51123),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__11771 (
            .O(N__51120),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    CascadeMux I__11770 (
            .O(N__51117),
            .I(N__51112));
    InMux I__11769 (
            .O(N__51116),
            .I(N__51109));
    InMux I__11768 (
            .O(N__51115),
            .I(N__51106));
    InMux I__11767 (
            .O(N__51112),
            .I(N__51103));
    LocalMux I__11766 (
            .O(N__51109),
            .I(N__51100));
    LocalMux I__11765 (
            .O(N__51106),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__11764 (
            .O(N__51103),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    Odrv12 I__11763 (
            .O(N__51100),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__11762 (
            .O(N__51093),
            .I(N__51090));
    LocalMux I__11761 (
            .O(N__51090),
            .I(N__51087));
    Odrv12 I__11760 (
            .O(N__51087),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__11759 (
            .O(N__51084),
            .I(bfn_20_27_0_));
    InMux I__11758 (
            .O(N__51081),
            .I(N__51077));
    InMux I__11757 (
            .O(N__51080),
            .I(N__51074));
    LocalMux I__11756 (
            .O(N__51077),
            .I(N__51071));
    LocalMux I__11755 (
            .O(N__51074),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv12 I__11754 (
            .O(N__51071),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__11753 (
            .O(N__51066),
            .I(N__51063));
    LocalMux I__11752 (
            .O(N__51063),
            .I(N__51060));
    Span4Mux_h I__11751 (
            .O(N__51060),
            .I(N__51057));
    Odrv4 I__11750 (
            .O(N__51057),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__11749 (
            .O(N__51054),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__11748 (
            .O(N__51051),
            .I(N__51048));
    LocalMux I__11747 (
            .O(N__51048),
            .I(N__51045));
    Span4Mux_v I__11746 (
            .O(N__51045),
            .I(N__51042));
    Span4Mux_h I__11745 (
            .O(N__51042),
            .I(N__51039));
    Odrv4 I__11744 (
            .O(N__51039),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__11743 (
            .O(N__51036),
            .I(N__51033));
    LocalMux I__11742 (
            .O(N__51033),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__11741 (
            .O(N__51030),
            .I(N__51027));
    LocalMux I__11740 (
            .O(N__51027),
            .I(N__51024));
    Span4Mux_v I__11739 (
            .O(N__51024),
            .I(N__51021));
    Span4Mux_h I__11738 (
            .O(N__51021),
            .I(N__51018));
    Odrv4 I__11737 (
            .O(N__51018),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__11736 (
            .O(N__51015),
            .I(N__51012));
    LocalMux I__11735 (
            .O(N__51012),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__11734 (
            .O(N__51009),
            .I(N__51006));
    LocalMux I__11733 (
            .O(N__51006),
            .I(N__51003));
    Span4Mux_h I__11732 (
            .O(N__51003),
            .I(N__51000));
    Span4Mux_h I__11731 (
            .O(N__51000),
            .I(N__50997));
    Odrv4 I__11730 (
            .O(N__50997),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__11729 (
            .O(N__50994),
            .I(N__50991));
    LocalMux I__11728 (
            .O(N__50991),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__11727 (
            .O(N__50988),
            .I(N__50985));
    LocalMux I__11726 (
            .O(N__50985),
            .I(N__50982));
    Span4Mux_h I__11725 (
            .O(N__50982),
            .I(N__50979));
    Span4Mux_h I__11724 (
            .O(N__50979),
            .I(N__50976));
    Odrv4 I__11723 (
            .O(N__50976),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__11722 (
            .O(N__50973),
            .I(N__50970));
    LocalMux I__11721 (
            .O(N__50970),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__11720 (
            .O(N__50967),
            .I(N__50964));
    LocalMux I__11719 (
            .O(N__50964),
            .I(N__50961));
    Span4Mux_v I__11718 (
            .O(N__50961),
            .I(N__50958));
    Span4Mux_h I__11717 (
            .O(N__50958),
            .I(N__50955));
    Odrv4 I__11716 (
            .O(N__50955),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__11715 (
            .O(N__50952),
            .I(N__50949));
    LocalMux I__11714 (
            .O(N__50949),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__11713 (
            .O(N__50946),
            .I(N__50943));
    LocalMux I__11712 (
            .O(N__50943),
            .I(N__50940));
    Span4Mux_h I__11711 (
            .O(N__50940),
            .I(N__50937));
    Span4Mux_h I__11710 (
            .O(N__50937),
            .I(N__50934));
    Odrv4 I__11709 (
            .O(N__50934),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__11708 (
            .O(N__50931),
            .I(N__50928));
    LocalMux I__11707 (
            .O(N__50928),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__11706 (
            .O(N__50925),
            .I(N__50922));
    LocalMux I__11705 (
            .O(N__50922),
            .I(N__50919));
    Span12Mux_s6_v I__11704 (
            .O(N__50919),
            .I(N__50916));
    Odrv12 I__11703 (
            .O(N__50916),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__11702 (
            .O(N__50913),
            .I(N__50910));
    LocalMux I__11701 (
            .O(N__50910),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__11700 (
            .O(N__50907),
            .I(N__50904));
    LocalMux I__11699 (
            .O(N__50904),
            .I(N__50901));
    Odrv4 I__11698 (
            .O(N__50901),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    InMux I__11697 (
            .O(N__50898),
            .I(N__50895));
    LocalMux I__11696 (
            .O(N__50895),
            .I(N__50892));
    Span4Mux_h I__11695 (
            .O(N__50892),
            .I(N__50888));
    InMux I__11694 (
            .O(N__50891),
            .I(N__50885));
    Odrv4 I__11693 (
            .O(N__50888),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__11692 (
            .O(N__50885),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    CascadeMux I__11691 (
            .O(N__50880),
            .I(N__50870));
    InMux I__11690 (
            .O(N__50879),
            .I(N__50866));
    InMux I__11689 (
            .O(N__50878),
            .I(N__50861));
    InMux I__11688 (
            .O(N__50877),
            .I(N__50861));
    InMux I__11687 (
            .O(N__50876),
            .I(N__50856));
    InMux I__11686 (
            .O(N__50875),
            .I(N__50856));
    InMux I__11685 (
            .O(N__50874),
            .I(N__50853));
    InMux I__11684 (
            .O(N__50873),
            .I(N__50838));
    InMux I__11683 (
            .O(N__50870),
            .I(N__50838));
    InMux I__11682 (
            .O(N__50869),
            .I(N__50838));
    LocalMux I__11681 (
            .O(N__50866),
            .I(N__50826));
    LocalMux I__11680 (
            .O(N__50861),
            .I(N__50826));
    LocalMux I__11679 (
            .O(N__50856),
            .I(N__50826));
    LocalMux I__11678 (
            .O(N__50853),
            .I(N__50819));
    InMux I__11677 (
            .O(N__50852),
            .I(N__50804));
    InMux I__11676 (
            .O(N__50851),
            .I(N__50804));
    InMux I__11675 (
            .O(N__50850),
            .I(N__50804));
    InMux I__11674 (
            .O(N__50849),
            .I(N__50804));
    InMux I__11673 (
            .O(N__50848),
            .I(N__50804));
    InMux I__11672 (
            .O(N__50847),
            .I(N__50799));
    InMux I__11671 (
            .O(N__50846),
            .I(N__50799));
    InMux I__11670 (
            .O(N__50845),
            .I(N__50796));
    LocalMux I__11669 (
            .O(N__50838),
            .I(N__50793));
    InMux I__11668 (
            .O(N__50837),
            .I(N__50788));
    InMux I__11667 (
            .O(N__50836),
            .I(N__50788));
    InMux I__11666 (
            .O(N__50835),
            .I(N__50785));
    InMux I__11665 (
            .O(N__50834),
            .I(N__50780));
    InMux I__11664 (
            .O(N__50833),
            .I(N__50780));
    Span4Mux_v I__11663 (
            .O(N__50826),
            .I(N__50777));
    InMux I__11662 (
            .O(N__50825),
            .I(N__50768));
    InMux I__11661 (
            .O(N__50824),
            .I(N__50768));
    InMux I__11660 (
            .O(N__50823),
            .I(N__50768));
    InMux I__11659 (
            .O(N__50822),
            .I(N__50768));
    Span4Mux_h I__11658 (
            .O(N__50819),
            .I(N__50765));
    InMux I__11657 (
            .O(N__50818),
            .I(N__50756));
    InMux I__11656 (
            .O(N__50817),
            .I(N__50756));
    InMux I__11655 (
            .O(N__50816),
            .I(N__50756));
    InMux I__11654 (
            .O(N__50815),
            .I(N__50756));
    LocalMux I__11653 (
            .O(N__50804),
            .I(N__50751));
    LocalMux I__11652 (
            .O(N__50799),
            .I(N__50751));
    LocalMux I__11651 (
            .O(N__50796),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11650 (
            .O(N__50793),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11649 (
            .O(N__50788),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11648 (
            .O(N__50785),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11647 (
            .O(N__50780),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11646 (
            .O(N__50777),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11645 (
            .O(N__50768),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11644 (
            .O(N__50765),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11643 (
            .O(N__50756),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11642 (
            .O(N__50751),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__11641 (
            .O(N__50730),
            .I(N__50727));
    LocalMux I__11640 (
            .O(N__50727),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    CascadeMux I__11639 (
            .O(N__50724),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_));
    InMux I__11638 (
            .O(N__50721),
            .I(N__50718));
    LocalMux I__11637 (
            .O(N__50718),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ));
    InMux I__11636 (
            .O(N__50715),
            .I(N__50712));
    LocalMux I__11635 (
            .O(N__50712),
            .I(N__50709));
    Span4Mux_h I__11634 (
            .O(N__50709),
            .I(N__50705));
    InMux I__11633 (
            .O(N__50708),
            .I(N__50702));
    Odrv4 I__11632 (
            .O(N__50705),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__11631 (
            .O(N__50702),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__11630 (
            .O(N__50697),
            .I(N__50693));
    CascadeMux I__11629 (
            .O(N__50696),
            .I(N__50690));
    LocalMux I__11628 (
            .O(N__50693),
            .I(N__50687));
    InMux I__11627 (
            .O(N__50690),
            .I(N__50684));
    Odrv4 I__11626 (
            .O(N__50687),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__11625 (
            .O(N__50684),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__11624 (
            .O(N__50679),
            .I(N__50676));
    LocalMux I__11623 (
            .O(N__50676),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ));
    CascadeMux I__11622 (
            .O(N__50673),
            .I(N__50669));
    InMux I__11621 (
            .O(N__50672),
            .I(N__50666));
    InMux I__11620 (
            .O(N__50669),
            .I(N__50663));
    LocalMux I__11619 (
            .O(N__50666),
            .I(N__50657));
    LocalMux I__11618 (
            .O(N__50663),
            .I(N__50657));
    InMux I__11617 (
            .O(N__50662),
            .I(N__50654));
    Span4Mux_h I__11616 (
            .O(N__50657),
            .I(N__50651));
    LocalMux I__11615 (
            .O(N__50654),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__11614 (
            .O(N__50651),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__11613 (
            .O(N__50646),
            .I(N__50643));
    LocalMux I__11612 (
            .O(N__50643),
            .I(N__50640));
    Span4Mux_h I__11611 (
            .O(N__50640),
            .I(N__50636));
    InMux I__11610 (
            .O(N__50639),
            .I(N__50633));
    Odrv4 I__11609 (
            .O(N__50636),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__11608 (
            .O(N__50633),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CascadeMux I__11607 (
            .O(N__50628),
            .I(N__50624));
    InMux I__11606 (
            .O(N__50627),
            .I(N__50621));
    InMux I__11605 (
            .O(N__50624),
            .I(N__50618));
    LocalMux I__11604 (
            .O(N__50621),
            .I(N__50612));
    LocalMux I__11603 (
            .O(N__50618),
            .I(N__50612));
    InMux I__11602 (
            .O(N__50617),
            .I(N__50609));
    Span4Mux_h I__11601 (
            .O(N__50612),
            .I(N__50606));
    LocalMux I__11600 (
            .O(N__50609),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__11599 (
            .O(N__50606),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__11598 (
            .O(N__50601),
            .I(N__50598));
    LocalMux I__11597 (
            .O(N__50598),
            .I(N__50595));
    Span4Mux_v I__11596 (
            .O(N__50595),
            .I(N__50591));
    InMux I__11595 (
            .O(N__50594),
            .I(N__50588));
    Odrv4 I__11594 (
            .O(N__50591),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__11593 (
            .O(N__50588),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    CEMux I__11592 (
            .O(N__50583),
            .I(N__50579));
    CEMux I__11591 (
            .O(N__50582),
            .I(N__50576));
    LocalMux I__11590 (
            .O(N__50579),
            .I(N__50570));
    LocalMux I__11589 (
            .O(N__50576),
            .I(N__50567));
    CEMux I__11588 (
            .O(N__50575),
            .I(N__50564));
    CEMux I__11587 (
            .O(N__50574),
            .I(N__50561));
    CEMux I__11586 (
            .O(N__50573),
            .I(N__50558));
    Span4Mux_h I__11585 (
            .O(N__50570),
            .I(N__50549));
    Span4Mux_v I__11584 (
            .O(N__50567),
            .I(N__50549));
    LocalMux I__11583 (
            .O(N__50564),
            .I(N__50549));
    LocalMux I__11582 (
            .O(N__50561),
            .I(N__50549));
    LocalMux I__11581 (
            .O(N__50558),
            .I(N__50546));
    Odrv4 I__11580 (
            .O(N__50549),
            .I(\delay_measurement_inst.delay_hc_timer.N_155_i ));
    Odrv4 I__11579 (
            .O(N__50546),
            .I(\delay_measurement_inst.delay_hc_timer.N_155_i ));
    InMux I__11578 (
            .O(N__50541),
            .I(N__50538));
    LocalMux I__11577 (
            .O(N__50538),
            .I(N__50535));
    Span4Mux_v I__11576 (
            .O(N__50535),
            .I(N__50532));
    Span4Mux_h I__11575 (
            .O(N__50532),
            .I(N__50529));
    Odrv4 I__11574 (
            .O(N__50529),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__11573 (
            .O(N__50526),
            .I(N__50523));
    LocalMux I__11572 (
            .O(N__50523),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__11571 (
            .O(N__50520),
            .I(N__50517));
    LocalMux I__11570 (
            .O(N__50517),
            .I(N__50514));
    Span12Mux_s7_v I__11569 (
            .O(N__50514),
            .I(N__50511));
    Odrv12 I__11568 (
            .O(N__50511),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__11567 (
            .O(N__50508),
            .I(N__50505));
    LocalMux I__11566 (
            .O(N__50505),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__11565 (
            .O(N__50502),
            .I(N__50499));
    LocalMux I__11564 (
            .O(N__50499),
            .I(N__50496));
    Span12Mux_h I__11563 (
            .O(N__50496),
            .I(N__50493));
    Odrv12 I__11562 (
            .O(N__50493),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__11561 (
            .O(N__50490),
            .I(N__50487));
    LocalMux I__11560 (
            .O(N__50487),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__11559 (
            .O(N__50484),
            .I(N__50481));
    LocalMux I__11558 (
            .O(N__50481),
            .I(N__50478));
    Span4Mux_v I__11557 (
            .O(N__50478),
            .I(N__50474));
    InMux I__11556 (
            .O(N__50477),
            .I(N__50471));
    Odrv4 I__11555 (
            .O(N__50474),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__11554 (
            .O(N__50471),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__11553 (
            .O(N__50466),
            .I(N__50463));
    LocalMux I__11552 (
            .O(N__50463),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    CascadeMux I__11551 (
            .O(N__50460),
            .I(elapsed_time_ns_1_RNI14DN9_0_23_cascade_));
    InMux I__11550 (
            .O(N__50457),
            .I(N__50454));
    LocalMux I__11549 (
            .O(N__50454),
            .I(N__50451));
    Odrv4 I__11548 (
            .O(N__50451),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ));
    InMux I__11547 (
            .O(N__50448),
            .I(N__50444));
    InMux I__11546 (
            .O(N__50447),
            .I(N__50441));
    LocalMux I__11545 (
            .O(N__50444),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__11544 (
            .O(N__50441),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__11543 (
            .O(N__50436),
            .I(N__50433));
    LocalMux I__11542 (
            .O(N__50433),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ));
    InMux I__11541 (
            .O(N__50430),
            .I(N__50427));
    LocalMux I__11540 (
            .O(N__50427),
            .I(N__50423));
    InMux I__11539 (
            .O(N__50426),
            .I(N__50420));
    Odrv4 I__11538 (
            .O(N__50423),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__11537 (
            .O(N__50420),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__11536 (
            .O(N__50415),
            .I(N__50411));
    InMux I__11535 (
            .O(N__50414),
            .I(N__50408));
    LocalMux I__11534 (
            .O(N__50411),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__11533 (
            .O(N__50408),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__11532 (
            .O(N__50403),
            .I(N__50400));
    LocalMux I__11531 (
            .O(N__50400),
            .I(N__50397));
    Span4Mux_v I__11530 (
            .O(N__50397),
            .I(N__50393));
    InMux I__11529 (
            .O(N__50396),
            .I(N__50390));
    Odrv4 I__11528 (
            .O(N__50393),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__11527 (
            .O(N__50390),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__11526 (
            .O(N__50385),
            .I(N__50382));
    LocalMux I__11525 (
            .O(N__50382),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    CascadeMux I__11524 (
            .O(N__50379),
            .I(elapsed_time_ns_1_RNI58DN9_0_27_cascade_));
    InMux I__11523 (
            .O(N__50376),
            .I(N__50373));
    LocalMux I__11522 (
            .O(N__50373),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ));
    InMux I__11521 (
            .O(N__50370),
            .I(N__50366));
    InMux I__11520 (
            .O(N__50369),
            .I(N__50363));
    LocalMux I__11519 (
            .O(N__50366),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__11518 (
            .O(N__50363),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__11517 (
            .O(N__50358),
            .I(N__50355));
    LocalMux I__11516 (
            .O(N__50355),
            .I(N__50351));
    InMux I__11515 (
            .O(N__50354),
            .I(N__50348));
    Odrv4 I__11514 (
            .O(N__50351),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__11513 (
            .O(N__50348),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__11512 (
            .O(N__50343),
            .I(N__50340));
    LocalMux I__11511 (
            .O(N__50340),
            .I(N__50337));
    Span4Mux_h I__11510 (
            .O(N__50337),
            .I(N__50333));
    InMux I__11509 (
            .O(N__50336),
            .I(N__50330));
    Odrv4 I__11508 (
            .O(N__50333),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__11507 (
            .O(N__50330),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__11506 (
            .O(N__50325),
            .I(N__50322));
    LocalMux I__11505 (
            .O(N__50322),
            .I(N__50318));
    InMux I__11504 (
            .O(N__50321),
            .I(N__50315));
    Odrv4 I__11503 (
            .O(N__50318),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__11502 (
            .O(N__50315),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    CascadeMux I__11501 (
            .O(N__50310),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ));
    InMux I__11500 (
            .O(N__50307),
            .I(N__50300));
    InMux I__11499 (
            .O(N__50306),
            .I(N__50300));
    InMux I__11498 (
            .O(N__50305),
            .I(N__50297));
    LocalMux I__11497 (
            .O(N__50300),
            .I(N__50294));
    LocalMux I__11496 (
            .O(N__50297),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ));
    Odrv12 I__11495 (
            .O(N__50294),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ));
    CascadeMux I__11494 (
            .O(N__50289),
            .I(N__50285));
    CascadeMux I__11493 (
            .O(N__50288),
            .I(N__50282));
    InMux I__11492 (
            .O(N__50285),
            .I(N__50277));
    InMux I__11491 (
            .O(N__50282),
            .I(N__50277));
    LocalMux I__11490 (
            .O(N__50277),
            .I(N__50273));
    InMux I__11489 (
            .O(N__50276),
            .I(N__50270));
    Span4Mux_h I__11488 (
            .O(N__50273),
            .I(N__50267));
    LocalMux I__11487 (
            .O(N__50270),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ));
    Odrv4 I__11486 (
            .O(N__50267),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ));
    CascadeMux I__11485 (
            .O(N__50262),
            .I(N__50259));
    InMux I__11484 (
            .O(N__50259),
            .I(N__50256));
    LocalMux I__11483 (
            .O(N__50256),
            .I(N__50253));
    Span4Mux_h I__11482 (
            .O(N__50253),
            .I(N__50250));
    Odrv4 I__11481 (
            .O(N__50250),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ));
    InMux I__11480 (
            .O(N__50247),
            .I(N__50243));
    InMux I__11479 (
            .O(N__50246),
            .I(N__50240));
    LocalMux I__11478 (
            .O(N__50243),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_27));
    LocalMux I__11477 (
            .O(N__50240),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_27));
    InMux I__11476 (
            .O(N__50235),
            .I(N__50229));
    InMux I__11475 (
            .O(N__50234),
            .I(N__50229));
    LocalMux I__11474 (
            .O(N__50229),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ));
    InMux I__11473 (
            .O(N__50226),
            .I(N__50222));
    InMux I__11472 (
            .O(N__50225),
            .I(N__50219));
    LocalMux I__11471 (
            .O(N__50222),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_26));
    LocalMux I__11470 (
            .O(N__50219),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_26));
    InMux I__11469 (
            .O(N__50214),
            .I(N__50208));
    InMux I__11468 (
            .O(N__50213),
            .I(N__50208));
    LocalMux I__11467 (
            .O(N__50208),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ));
    InMux I__11466 (
            .O(N__50205),
            .I(N__50201));
    InMux I__11465 (
            .O(N__50204),
            .I(N__50198));
    LocalMux I__11464 (
            .O(N__50201),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_24));
    LocalMux I__11463 (
            .O(N__50198),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_24));
    InMux I__11462 (
            .O(N__50193),
            .I(N__50187));
    InMux I__11461 (
            .O(N__50192),
            .I(N__50187));
    LocalMux I__11460 (
            .O(N__50187),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ));
    InMux I__11459 (
            .O(N__50184),
            .I(N__50180));
    InMux I__11458 (
            .O(N__50183),
            .I(N__50177));
    LocalMux I__11457 (
            .O(N__50180),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_25));
    LocalMux I__11456 (
            .O(N__50177),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_25));
    CascadeMux I__11455 (
            .O(N__50172),
            .I(N__50168));
    CascadeMux I__11454 (
            .O(N__50171),
            .I(N__50165));
    InMux I__11453 (
            .O(N__50168),
            .I(N__50160));
    InMux I__11452 (
            .O(N__50165),
            .I(N__50160));
    LocalMux I__11451 (
            .O(N__50160),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ));
    CEMux I__11450 (
            .O(N__50157),
            .I(N__50152));
    CEMux I__11449 (
            .O(N__50156),
            .I(N__50149));
    CEMux I__11448 (
            .O(N__50155),
            .I(N__50142));
    LocalMux I__11447 (
            .O(N__50152),
            .I(N__50135));
    LocalMux I__11446 (
            .O(N__50149),
            .I(N__50135));
    CEMux I__11445 (
            .O(N__50148),
            .I(N__50132));
    CEMux I__11444 (
            .O(N__50147),
            .I(N__50128));
    CEMux I__11443 (
            .O(N__50146),
            .I(N__50125));
    CEMux I__11442 (
            .O(N__50145),
            .I(N__50122));
    LocalMux I__11441 (
            .O(N__50142),
            .I(N__50119));
    CEMux I__11440 (
            .O(N__50141),
            .I(N__50116));
    CEMux I__11439 (
            .O(N__50140),
            .I(N__50113));
    Span4Mux_v I__11438 (
            .O(N__50135),
            .I(N__50108));
    LocalMux I__11437 (
            .O(N__50132),
            .I(N__50108));
    CEMux I__11436 (
            .O(N__50131),
            .I(N__50105));
    LocalMux I__11435 (
            .O(N__50128),
            .I(N__50098));
    LocalMux I__11434 (
            .O(N__50125),
            .I(N__50098));
    LocalMux I__11433 (
            .O(N__50122),
            .I(N__50098));
    Span4Mux_v I__11432 (
            .O(N__50119),
            .I(N__50095));
    LocalMux I__11431 (
            .O(N__50116),
            .I(N__50088));
    LocalMux I__11430 (
            .O(N__50113),
            .I(N__50088));
    Span4Mux_v I__11429 (
            .O(N__50108),
            .I(N__50088));
    LocalMux I__11428 (
            .O(N__50105),
            .I(N__50085));
    Span4Mux_v I__11427 (
            .O(N__50098),
            .I(N__50082));
    Span4Mux_v I__11426 (
            .O(N__50095),
            .I(N__50077));
    Span4Mux_v I__11425 (
            .O(N__50088),
            .I(N__50077));
    Span12Mux_v I__11424 (
            .O(N__50085),
            .I(N__50074));
    Span4Mux_h I__11423 (
            .O(N__50082),
            .I(N__50071));
    Span4Mux_h I__11422 (
            .O(N__50077),
            .I(N__50068));
    Odrv12 I__11421 (
            .O(N__50074),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__11420 (
            .O(N__50071),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__11419 (
            .O(N__50068),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    InMux I__11418 (
            .O(N__50061),
            .I(N__50058));
    LocalMux I__11417 (
            .O(N__50058),
            .I(N__50054));
    CascadeMux I__11416 (
            .O(N__50057),
            .I(N__50051));
    Span4Mux_v I__11415 (
            .O(N__50054),
            .I(N__50048));
    InMux I__11414 (
            .O(N__50051),
            .I(N__50045));
    Odrv4 I__11413 (
            .O(N__50048),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__11412 (
            .O(N__50045),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__11411 (
            .O(N__50040),
            .I(N__50037));
    LocalMux I__11410 (
            .O(N__50037),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    CascadeMux I__11409 (
            .O(N__50034),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_));
    InMux I__11408 (
            .O(N__50031),
            .I(N__50028));
    LocalMux I__11407 (
            .O(N__50028),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ));
    InMux I__11406 (
            .O(N__50025),
            .I(N__50022));
    LocalMux I__11405 (
            .O(N__50022),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ));
    InMux I__11404 (
            .O(N__50019),
            .I(N__50016));
    LocalMux I__11403 (
            .O(N__50016),
            .I(N__50012));
    InMux I__11402 (
            .O(N__50015),
            .I(N__50009));
    Odrv4 I__11401 (
            .O(N__50012),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_19));
    LocalMux I__11400 (
            .O(N__50009),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_19));
    InMux I__11399 (
            .O(N__50004),
            .I(N__50001));
    LocalMux I__11398 (
            .O(N__50001),
            .I(N__49998));
    Span4Mux_h I__11397 (
            .O(N__49998),
            .I(N__49995));
    Odrv4 I__11396 (
            .O(N__49995),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt16 ));
    InMux I__11395 (
            .O(N__49992),
            .I(N__49986));
    InMux I__11394 (
            .O(N__49991),
            .I(N__49986));
    LocalMux I__11393 (
            .O(N__49986),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ));
    InMux I__11392 (
            .O(N__49983),
            .I(N__49976));
    InMux I__11391 (
            .O(N__49982),
            .I(N__49976));
    InMux I__11390 (
            .O(N__49981),
            .I(N__49973));
    LocalMux I__11389 (
            .O(N__49976),
            .I(N__49970));
    LocalMux I__11388 (
            .O(N__49973),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ));
    Odrv12 I__11387 (
            .O(N__49970),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ));
    CascadeMux I__11386 (
            .O(N__49965),
            .I(N__49961));
    CascadeMux I__11385 (
            .O(N__49964),
            .I(N__49958));
    InMux I__11384 (
            .O(N__49961),
            .I(N__49952));
    InMux I__11383 (
            .O(N__49958),
            .I(N__49952));
    InMux I__11382 (
            .O(N__49957),
            .I(N__49949));
    LocalMux I__11381 (
            .O(N__49952),
            .I(N__49946));
    LocalMux I__11380 (
            .O(N__49949),
            .I(N__49941));
    Span4Mux_h I__11379 (
            .O(N__49946),
            .I(N__49941));
    Odrv4 I__11378 (
            .O(N__49941),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ));
    CascadeMux I__11377 (
            .O(N__49938),
            .I(N__49935));
    InMux I__11376 (
            .O(N__49935),
            .I(N__49932));
    LocalMux I__11375 (
            .O(N__49932),
            .I(N__49929));
    Span4Mux_h I__11374 (
            .O(N__49929),
            .I(N__49926));
    Odrv4 I__11373 (
            .O(N__49926),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ));
    InMux I__11372 (
            .O(N__49923),
            .I(N__49920));
    LocalMux I__11371 (
            .O(N__49920),
            .I(N__49917));
    Span4Mux_v I__11370 (
            .O(N__49917),
            .I(N__49913));
    InMux I__11369 (
            .O(N__49916),
            .I(N__49910));
    Odrv4 I__11368 (
            .O(N__49913),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_17));
    LocalMux I__11367 (
            .O(N__49910),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_17));
    InMux I__11366 (
            .O(N__49905),
            .I(N__49899));
    InMux I__11365 (
            .O(N__49904),
            .I(N__49899));
    LocalMux I__11364 (
            .O(N__49899),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ));
    CascadeMux I__11363 (
            .O(N__49896),
            .I(N__49893));
    InMux I__11362 (
            .O(N__49893),
            .I(N__49890));
    LocalMux I__11361 (
            .O(N__49890),
            .I(N__49887));
    Span4Mux_v I__11360 (
            .O(N__49887),
            .I(N__49884));
    Odrv4 I__11359 (
            .O(N__49884),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt18 ));
    InMux I__11358 (
            .O(N__49881),
            .I(N__49875));
    InMux I__11357 (
            .O(N__49880),
            .I(N__49875));
    LocalMux I__11356 (
            .O(N__49875),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ));
    InMux I__11355 (
            .O(N__49872),
            .I(N__49866));
    InMux I__11354 (
            .O(N__49871),
            .I(N__49866));
    LocalMux I__11353 (
            .O(N__49866),
            .I(N__49862));
    InMux I__11352 (
            .O(N__49865),
            .I(N__49859));
    Span4Mux_h I__11351 (
            .O(N__49862),
            .I(N__49856));
    LocalMux I__11350 (
            .O(N__49859),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__11349 (
            .O(N__49856),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    CascadeMux I__11348 (
            .O(N__49851),
            .I(N__49847));
    CascadeMux I__11347 (
            .O(N__49850),
            .I(N__49844));
    InMux I__11346 (
            .O(N__49847),
            .I(N__49838));
    InMux I__11345 (
            .O(N__49844),
            .I(N__49838));
    InMux I__11344 (
            .O(N__49843),
            .I(N__49835));
    LocalMux I__11343 (
            .O(N__49838),
            .I(N__49832));
    LocalMux I__11342 (
            .O(N__49835),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    Odrv12 I__11341 (
            .O(N__49832),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    InMux I__11340 (
            .O(N__49827),
            .I(N__49821));
    InMux I__11339 (
            .O(N__49826),
            .I(N__49821));
    LocalMux I__11338 (
            .O(N__49821),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ));
    InMux I__11337 (
            .O(N__49818),
            .I(N__49815));
    LocalMux I__11336 (
            .O(N__49815),
            .I(N__49812));
    Span4Mux_h I__11335 (
            .O(N__49812),
            .I(N__49809));
    Odrv4 I__11334 (
            .O(N__49809),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ));
    CascadeMux I__11333 (
            .O(N__49806),
            .I(N__49803));
    InMux I__11332 (
            .O(N__49803),
            .I(N__49800));
    LocalMux I__11331 (
            .O(N__49800),
            .I(N__49797));
    Span4Mux_h I__11330 (
            .O(N__49797),
            .I(N__49794));
    Odrv4 I__11329 (
            .O(N__49794),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt24 ));
    InMux I__11328 (
            .O(N__49791),
            .I(N__49784));
    InMux I__11327 (
            .O(N__49790),
            .I(N__49784));
    InMux I__11326 (
            .O(N__49789),
            .I(N__49781));
    LocalMux I__11325 (
            .O(N__49784),
            .I(N__49778));
    LocalMux I__11324 (
            .O(N__49781),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ));
    Odrv12 I__11323 (
            .O(N__49778),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ));
    InMux I__11322 (
            .O(N__49773),
            .I(N__49766));
    InMux I__11321 (
            .O(N__49772),
            .I(N__49766));
    InMux I__11320 (
            .O(N__49771),
            .I(N__49763));
    LocalMux I__11319 (
            .O(N__49766),
            .I(N__49760));
    LocalMux I__11318 (
            .O(N__49763),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ));
    Odrv12 I__11317 (
            .O(N__49760),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ));
    InMux I__11316 (
            .O(N__49755),
            .I(N__49752));
    LocalMux I__11315 (
            .O(N__49752),
            .I(N__49749));
    Odrv12 I__11314 (
            .O(N__49749),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ));
    InMux I__11313 (
            .O(N__49746),
            .I(N__49743));
    LocalMux I__11312 (
            .O(N__49743),
            .I(N__49740));
    Odrv12 I__11311 (
            .O(N__49740),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt26 ));
    InMux I__11310 (
            .O(N__49737),
            .I(N__49734));
    LocalMux I__11309 (
            .O(N__49734),
            .I(\pwm_generator_inst.un19_threshold_0_axb_7 ));
    CascadeMux I__11308 (
            .O(N__49731),
            .I(N__49728));
    InMux I__11307 (
            .O(N__49728),
            .I(N__49725));
    LocalMux I__11306 (
            .O(N__49725),
            .I(N__49722));
    Span4Mux_v I__11305 (
            .O(N__49722),
            .I(N__49719));
    Odrv4 I__11304 (
            .O(N__49719),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__11303 (
            .O(N__49716),
            .I(\pwm_generator_inst.un19_threshold_0_cry_6 ));
    CascadeMux I__11302 (
            .O(N__49713),
            .I(N__49710));
    InMux I__11301 (
            .O(N__49710),
            .I(N__49707));
    LocalMux I__11300 (
            .O(N__49707),
            .I(N__49704));
    Odrv12 I__11299 (
            .O(N__49704),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__11298 (
            .O(N__49701),
            .I(bfn_17_27_0_));
    InMux I__11297 (
            .O(N__49698),
            .I(N__49695));
    LocalMux I__11296 (
            .O(N__49695),
            .I(N__49692));
    Span4Mux_h I__11295 (
            .O(N__49692),
            .I(N__49689));
    Odrv4 I__11294 (
            .O(N__49689),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__11293 (
            .O(N__49686),
            .I(\pwm_generator_inst.un19_threshold_0_cry_8 ));
    CascadeMux I__11292 (
            .O(N__49683),
            .I(N__49680));
    InMux I__11291 (
            .O(N__49680),
            .I(N__49677));
    LocalMux I__11290 (
            .O(N__49677),
            .I(N__49674));
    Odrv4 I__11289 (
            .O(N__49674),
            .I(\pwm_generator_inst.un14_counter_9 ));
    InMux I__11288 (
            .O(N__49671),
            .I(N__49668));
    LocalMux I__11287 (
            .O(N__49668),
            .I(N__49665));
    Span4Mux_h I__11286 (
            .O(N__49665),
            .I(N__49661));
    InMux I__11285 (
            .O(N__49664),
            .I(N__49658));
    Odrv4 I__11284 (
            .O(N__49661),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    LocalMux I__11283 (
            .O(N__49658),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__11282 (
            .O(N__49653),
            .I(N__49650));
    LocalMux I__11281 (
            .O(N__49650),
            .I(\pwm_generator_inst.un19_threshold_0_axb_6 ));
    CascadeMux I__11280 (
            .O(N__49647),
            .I(N__49644));
    InMux I__11279 (
            .O(N__49644),
            .I(N__49641));
    LocalMux I__11278 (
            .O(N__49641),
            .I(N__49637));
    InMux I__11277 (
            .O(N__49640),
            .I(N__49634));
    Span4Mux_h I__11276 (
            .O(N__49637),
            .I(N__49631));
    LocalMux I__11275 (
            .O(N__49634),
            .I(N__49628));
    Odrv4 I__11274 (
            .O(N__49631),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    Odrv4 I__11273 (
            .O(N__49628),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__11272 (
            .O(N__49623),
            .I(N__49620));
    LocalMux I__11271 (
            .O(N__49620),
            .I(\pwm_generator_inst.un19_threshold_0_axb_4 ));
    InMux I__11270 (
            .O(N__49617),
            .I(N__49614));
    LocalMux I__11269 (
            .O(N__49614),
            .I(N__49611));
    Span4Mux_h I__11268 (
            .O(N__49611),
            .I(N__49607));
    InMux I__11267 (
            .O(N__49610),
            .I(N__49604));
    Odrv4 I__11266 (
            .O(N__49607),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    LocalMux I__11265 (
            .O(N__49604),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    InMux I__11264 (
            .O(N__49599),
            .I(N__49596));
    LocalMux I__11263 (
            .O(N__49596),
            .I(\pwm_generator_inst.un19_threshold_0_axb_8 ));
    InMux I__11262 (
            .O(N__49593),
            .I(N__49590));
    LocalMux I__11261 (
            .O(N__49590),
            .I(N__49586));
    InMux I__11260 (
            .O(N__49589),
            .I(N__49583));
    Odrv4 I__11259 (
            .O(N__49586),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_16));
    LocalMux I__11258 (
            .O(N__49583),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_16));
    InMux I__11257 (
            .O(N__49578),
            .I(N__49574));
    InMux I__11256 (
            .O(N__49577),
            .I(N__49571));
    LocalMux I__11255 (
            .O(N__49574),
            .I(N__49568));
    LocalMux I__11254 (
            .O(N__49571),
            .I(N__49565));
    Span4Mux_h I__11253 (
            .O(N__49568),
            .I(N__49562));
    Odrv4 I__11252 (
            .O(N__49565),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_18));
    Odrv4 I__11251 (
            .O(N__49562),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_18));
    InMux I__11250 (
            .O(N__49557),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__11249 (
            .O(N__49554),
            .I(N__49551));
    LocalMux I__11248 (
            .O(N__49551),
            .I(N__49548));
    Span4Mux_s0_v I__11247 (
            .O(N__49548),
            .I(N__49545));
    Sp12to4 I__11246 (
            .O(N__49545),
            .I(N__49542));
    Span12Mux_h I__11245 (
            .O(N__49542),
            .I(N__49539));
    Span12Mux_v I__11244 (
            .O(N__49539),
            .I(N__49536));
    Span12Mux_v I__11243 (
            .O(N__49536),
            .I(N__49533));
    Odrv12 I__11242 (
            .O(N__49533),
            .I(pwm_output_c));
    InMux I__11241 (
            .O(N__49530),
            .I(N__49527));
    LocalMux I__11240 (
            .O(N__49527),
            .I(\pwm_generator_inst.un19_threshold_0_axb_0 ));
    CascadeMux I__11239 (
            .O(N__49524),
            .I(N__49521));
    InMux I__11238 (
            .O(N__49521),
            .I(N__49518));
    LocalMux I__11237 (
            .O(N__49518),
            .I(N__49515));
    Span4Mux_h I__11236 (
            .O(N__49515),
            .I(N__49512));
    Odrv4 I__11235 (
            .O(N__49512),
            .I(\pwm_generator_inst.un14_counter_0 ));
    CascadeMux I__11234 (
            .O(N__49509),
            .I(N__49506));
    InMux I__11233 (
            .O(N__49506),
            .I(N__49503));
    LocalMux I__11232 (
            .O(N__49503),
            .I(N__49500));
    Span4Mux_h I__11231 (
            .O(N__49500),
            .I(N__49497));
    Odrv4 I__11230 (
            .O(N__49497),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__11229 (
            .O(N__49494),
            .I(\pwm_generator_inst.un19_threshold_0_cry_0 ));
    CascadeMux I__11228 (
            .O(N__49491),
            .I(N__49488));
    InMux I__11227 (
            .O(N__49488),
            .I(N__49485));
    LocalMux I__11226 (
            .O(N__49485),
            .I(\pwm_generator_inst.un19_threshold_0_axb_2 ));
    CascadeMux I__11225 (
            .O(N__49482),
            .I(N__49479));
    InMux I__11224 (
            .O(N__49479),
            .I(N__49476));
    LocalMux I__11223 (
            .O(N__49476),
            .I(N__49473));
    Span4Mux_v I__11222 (
            .O(N__49473),
            .I(N__49470));
    Odrv4 I__11221 (
            .O(N__49470),
            .I(\pwm_generator_inst.un14_counter_2 ));
    InMux I__11220 (
            .O(N__49467),
            .I(\pwm_generator_inst.un19_threshold_0_cry_1 ));
    InMux I__11219 (
            .O(N__49464),
            .I(N__49461));
    LocalMux I__11218 (
            .O(N__49461),
            .I(\pwm_generator_inst.un19_threshold_0_axb_3 ));
    CascadeMux I__11217 (
            .O(N__49458),
            .I(N__49455));
    InMux I__11216 (
            .O(N__49455),
            .I(N__49452));
    LocalMux I__11215 (
            .O(N__49452),
            .I(N__49449));
    Span4Mux_v I__11214 (
            .O(N__49449),
            .I(N__49446));
    Odrv4 I__11213 (
            .O(N__49446),
            .I(\pwm_generator_inst.un14_counter_3 ));
    InMux I__11212 (
            .O(N__49443),
            .I(\pwm_generator_inst.un19_threshold_0_cry_2 ));
    CascadeMux I__11211 (
            .O(N__49440),
            .I(N__49437));
    InMux I__11210 (
            .O(N__49437),
            .I(N__49434));
    LocalMux I__11209 (
            .O(N__49434),
            .I(N__49431));
    Odrv4 I__11208 (
            .O(N__49431),
            .I(\pwm_generator_inst.un14_counter_4 ));
    InMux I__11207 (
            .O(N__49428),
            .I(\pwm_generator_inst.un19_threshold_0_cry_3 ));
    InMux I__11206 (
            .O(N__49425),
            .I(N__49422));
    LocalMux I__11205 (
            .O(N__49422),
            .I(\pwm_generator_inst.un19_threshold_0_axb_5 ));
    CascadeMux I__11204 (
            .O(N__49419),
            .I(N__49416));
    InMux I__11203 (
            .O(N__49416),
            .I(N__49413));
    LocalMux I__11202 (
            .O(N__49413),
            .I(N__49410));
    Span4Mux_v I__11201 (
            .O(N__49410),
            .I(N__49407));
    Odrv4 I__11200 (
            .O(N__49407),
            .I(\pwm_generator_inst.un14_counter_5 ));
    InMux I__11199 (
            .O(N__49404),
            .I(\pwm_generator_inst.un19_threshold_0_cry_4 ));
    CascadeMux I__11198 (
            .O(N__49401),
            .I(N__49398));
    InMux I__11197 (
            .O(N__49398),
            .I(N__49395));
    LocalMux I__11196 (
            .O(N__49395),
            .I(N__49392));
    Span4Mux_h I__11195 (
            .O(N__49392),
            .I(N__49389));
    Odrv4 I__11194 (
            .O(N__49389),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__11193 (
            .O(N__49386),
            .I(\pwm_generator_inst.un19_threshold_0_cry_5 ));
    InMux I__11192 (
            .O(N__49383),
            .I(N__49379));
    InMux I__11191 (
            .O(N__49382),
            .I(N__49375));
    LocalMux I__11190 (
            .O(N__49379),
            .I(N__49372));
    InMux I__11189 (
            .O(N__49378),
            .I(N__49369));
    LocalMux I__11188 (
            .O(N__49375),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__11187 (
            .O(N__49372),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__11186 (
            .O(N__49369),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__11185 (
            .O(N__49362),
            .I(N__49359));
    LocalMux I__11184 (
            .O(N__49359),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__11183 (
            .O(N__49356),
            .I(N__49352));
    InMux I__11182 (
            .O(N__49355),
            .I(N__49348));
    LocalMux I__11181 (
            .O(N__49352),
            .I(N__49345));
    InMux I__11180 (
            .O(N__49351),
            .I(N__49342));
    LocalMux I__11179 (
            .O(N__49348),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__11178 (
            .O(N__49345),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__11177 (
            .O(N__49342),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__11176 (
            .O(N__49335),
            .I(N__49332));
    LocalMux I__11175 (
            .O(N__49332),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__11174 (
            .O(N__49329),
            .I(N__49325));
    InMux I__11173 (
            .O(N__49328),
            .I(N__49321));
    LocalMux I__11172 (
            .O(N__49325),
            .I(N__49318));
    InMux I__11171 (
            .O(N__49324),
            .I(N__49315));
    LocalMux I__11170 (
            .O(N__49321),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__11169 (
            .O(N__49318),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__11168 (
            .O(N__49315),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__11167 (
            .O(N__49308),
            .I(N__49305));
    LocalMux I__11166 (
            .O(N__49305),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__11165 (
            .O(N__49302),
            .I(N__49298));
    InMux I__11164 (
            .O(N__49301),
            .I(N__49294));
    LocalMux I__11163 (
            .O(N__49298),
            .I(N__49291));
    InMux I__11162 (
            .O(N__49297),
            .I(N__49288));
    LocalMux I__11161 (
            .O(N__49294),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__11160 (
            .O(N__49291),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__11159 (
            .O(N__49288),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__11158 (
            .O(N__49281),
            .I(N__49278));
    LocalMux I__11157 (
            .O(N__49278),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__11156 (
            .O(N__49275),
            .I(N__49272));
    LocalMux I__11155 (
            .O(N__49272),
            .I(N__49267));
    InMux I__11154 (
            .O(N__49271),
            .I(N__49264));
    InMux I__11153 (
            .O(N__49270),
            .I(N__49261));
    Odrv4 I__11152 (
            .O(N__49267),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__11151 (
            .O(N__49264),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__11150 (
            .O(N__49261),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__11149 (
            .O(N__49254),
            .I(N__49251));
    LocalMux I__11148 (
            .O(N__49251),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__11147 (
            .O(N__49248),
            .I(N__49244));
    InMux I__11146 (
            .O(N__49247),
            .I(N__49240));
    LocalMux I__11145 (
            .O(N__49244),
            .I(N__49237));
    InMux I__11144 (
            .O(N__49243),
            .I(N__49234));
    LocalMux I__11143 (
            .O(N__49240),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__11142 (
            .O(N__49237),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__11141 (
            .O(N__49234),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__11140 (
            .O(N__49227),
            .I(N__49224));
    LocalMux I__11139 (
            .O(N__49224),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__11138 (
            .O(N__49221),
            .I(N__49216));
    InMux I__11137 (
            .O(N__49220),
            .I(N__49213));
    InMux I__11136 (
            .O(N__49219),
            .I(N__49210));
    LocalMux I__11135 (
            .O(N__49216),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__11134 (
            .O(N__49213),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__11133 (
            .O(N__49210),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__11132 (
            .O(N__49203),
            .I(N__49200));
    LocalMux I__11131 (
            .O(N__49200),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__11130 (
            .O(N__49197),
            .I(N__49192));
    InMux I__11129 (
            .O(N__49196),
            .I(N__49189));
    InMux I__11128 (
            .O(N__49195),
            .I(N__49186));
    LocalMux I__11127 (
            .O(N__49192),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__11126 (
            .O(N__49189),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__11125 (
            .O(N__49186),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__11124 (
            .O(N__49179),
            .I(N__49176));
    LocalMux I__11123 (
            .O(N__49176),
            .I(\pwm_generator_inst.counter_i_9 ));
    CascadeMux I__11122 (
            .O(N__49173),
            .I(N__49170));
    InMux I__11121 (
            .O(N__49170),
            .I(N__49167));
    LocalMux I__11120 (
            .O(N__49167),
            .I(N__49162));
    InMux I__11119 (
            .O(N__49166),
            .I(N__49159));
    InMux I__11118 (
            .O(N__49165),
            .I(N__49156));
    Span4Mux_h I__11117 (
            .O(N__49162),
            .I(N__49153));
    LocalMux I__11116 (
            .O(N__49159),
            .I(N__49150));
    LocalMux I__11115 (
            .O(N__49156),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__11114 (
            .O(N__49153),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv12 I__11113 (
            .O(N__49150),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__11112 (
            .O(N__49143),
            .I(bfn_17_23_0_));
    CascadeMux I__11111 (
            .O(N__49140),
            .I(N__49137));
    InMux I__11110 (
            .O(N__49137),
            .I(N__49133));
    CascadeMux I__11109 (
            .O(N__49136),
            .I(N__49130));
    LocalMux I__11108 (
            .O(N__49133),
            .I(N__49126));
    InMux I__11107 (
            .O(N__49130),
            .I(N__49123));
    InMux I__11106 (
            .O(N__49129),
            .I(N__49120));
    Span4Mux_h I__11105 (
            .O(N__49126),
            .I(N__49117));
    LocalMux I__11104 (
            .O(N__49123),
            .I(N__49114));
    LocalMux I__11103 (
            .O(N__49120),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__11102 (
            .O(N__49117),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv12 I__11101 (
            .O(N__49114),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__11100 (
            .O(N__49107),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__11099 (
            .O(N__49104),
            .I(N__49097));
    InMux I__11098 (
            .O(N__49103),
            .I(N__49097));
    InMux I__11097 (
            .O(N__49102),
            .I(N__49094));
    LocalMux I__11096 (
            .O(N__49097),
            .I(N__49091));
    LocalMux I__11095 (
            .O(N__49094),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv12 I__11094 (
            .O(N__49091),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__11093 (
            .O(N__49086),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__11092 (
            .O(N__49083),
            .I(N__49076));
    InMux I__11091 (
            .O(N__49082),
            .I(N__49076));
    InMux I__11090 (
            .O(N__49081),
            .I(N__49073));
    LocalMux I__11089 (
            .O(N__49076),
            .I(N__49070));
    LocalMux I__11088 (
            .O(N__49073),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__11087 (
            .O(N__49070),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__11086 (
            .O(N__49065),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    CascadeMux I__11085 (
            .O(N__49062),
            .I(N__49059));
    InMux I__11084 (
            .O(N__49059),
            .I(N__49055));
    InMux I__11083 (
            .O(N__49058),
            .I(N__49052));
    LocalMux I__11082 (
            .O(N__49055),
            .I(N__49049));
    LocalMux I__11081 (
            .O(N__49052),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv12 I__11080 (
            .O(N__49049),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__11079 (
            .O(N__49044),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__11078 (
            .O(N__49041),
            .I(N__49003));
    InMux I__11077 (
            .O(N__49040),
            .I(N__49003));
    InMux I__11076 (
            .O(N__49039),
            .I(N__49003));
    InMux I__11075 (
            .O(N__49038),
            .I(N__49003));
    InMux I__11074 (
            .O(N__49037),
            .I(N__48994));
    InMux I__11073 (
            .O(N__49036),
            .I(N__48994));
    InMux I__11072 (
            .O(N__49035),
            .I(N__48994));
    InMux I__11071 (
            .O(N__49034),
            .I(N__48994));
    InMux I__11070 (
            .O(N__49033),
            .I(N__48985));
    InMux I__11069 (
            .O(N__49032),
            .I(N__48985));
    InMux I__11068 (
            .O(N__49031),
            .I(N__48985));
    InMux I__11067 (
            .O(N__49030),
            .I(N__48985));
    InMux I__11066 (
            .O(N__49029),
            .I(N__48976));
    InMux I__11065 (
            .O(N__49028),
            .I(N__48976));
    InMux I__11064 (
            .O(N__49027),
            .I(N__48976));
    InMux I__11063 (
            .O(N__49026),
            .I(N__48976));
    InMux I__11062 (
            .O(N__49025),
            .I(N__48971));
    InMux I__11061 (
            .O(N__49024),
            .I(N__48971));
    InMux I__11060 (
            .O(N__49023),
            .I(N__48962));
    InMux I__11059 (
            .O(N__49022),
            .I(N__48962));
    InMux I__11058 (
            .O(N__49021),
            .I(N__48962));
    InMux I__11057 (
            .O(N__49020),
            .I(N__48962));
    InMux I__11056 (
            .O(N__49019),
            .I(N__48953));
    InMux I__11055 (
            .O(N__49018),
            .I(N__48953));
    InMux I__11054 (
            .O(N__49017),
            .I(N__48953));
    InMux I__11053 (
            .O(N__49016),
            .I(N__48953));
    InMux I__11052 (
            .O(N__49015),
            .I(N__48944));
    InMux I__11051 (
            .O(N__49014),
            .I(N__48944));
    InMux I__11050 (
            .O(N__49013),
            .I(N__48944));
    InMux I__11049 (
            .O(N__49012),
            .I(N__48944));
    LocalMux I__11048 (
            .O(N__49003),
            .I(N__48937));
    LocalMux I__11047 (
            .O(N__48994),
            .I(N__48937));
    LocalMux I__11046 (
            .O(N__48985),
            .I(N__48937));
    LocalMux I__11045 (
            .O(N__48976),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__11044 (
            .O(N__48971),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__11043 (
            .O(N__48962),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__11042 (
            .O(N__48953),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__11041 (
            .O(N__48944),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__11040 (
            .O(N__48937),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__11039 (
            .O(N__48924),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CascadeMux I__11038 (
            .O(N__48921),
            .I(N__48918));
    InMux I__11037 (
            .O(N__48918),
            .I(N__48914));
    InMux I__11036 (
            .O(N__48917),
            .I(N__48911));
    LocalMux I__11035 (
            .O(N__48914),
            .I(N__48908));
    LocalMux I__11034 (
            .O(N__48911),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv12 I__11033 (
            .O(N__48908),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CEMux I__11032 (
            .O(N__48903),
            .I(N__48899));
    CEMux I__11031 (
            .O(N__48902),
            .I(N__48895));
    LocalMux I__11030 (
            .O(N__48899),
            .I(N__48892));
    CEMux I__11029 (
            .O(N__48898),
            .I(N__48889));
    LocalMux I__11028 (
            .O(N__48895),
            .I(N__48885));
    Span4Mux_v I__11027 (
            .O(N__48892),
            .I(N__48882));
    LocalMux I__11026 (
            .O(N__48889),
            .I(N__48879));
    CEMux I__11025 (
            .O(N__48888),
            .I(N__48876));
    Span4Mux_h I__11024 (
            .O(N__48885),
            .I(N__48873));
    Span4Mux_h I__11023 (
            .O(N__48882),
            .I(N__48870));
    Span4Mux_h I__11022 (
            .O(N__48879),
            .I(N__48867));
    LocalMux I__11021 (
            .O(N__48876),
            .I(N__48864));
    Odrv4 I__11020 (
            .O(N__48873),
            .I(\delay_measurement_inst.delay_hc_timer.N_156_i ));
    Odrv4 I__11019 (
            .O(N__48870),
            .I(\delay_measurement_inst.delay_hc_timer.N_156_i ));
    Odrv4 I__11018 (
            .O(N__48867),
            .I(\delay_measurement_inst.delay_hc_timer.N_156_i ));
    Odrv12 I__11017 (
            .O(N__48864),
            .I(\delay_measurement_inst.delay_hc_timer.N_156_i ));
    InMux I__11016 (
            .O(N__48855),
            .I(N__48850));
    InMux I__11015 (
            .O(N__48854),
            .I(N__48847));
    InMux I__11014 (
            .O(N__48853),
            .I(N__48844));
    LocalMux I__11013 (
            .O(N__48850),
            .I(N__48841));
    LocalMux I__11012 (
            .O(N__48847),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__11011 (
            .O(N__48844),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__11010 (
            .O(N__48841),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__11009 (
            .O(N__48834),
            .I(N__48831));
    LocalMux I__11008 (
            .O(N__48831),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__11007 (
            .O(N__48828),
            .I(N__48823));
    InMux I__11006 (
            .O(N__48827),
            .I(N__48820));
    InMux I__11005 (
            .O(N__48826),
            .I(N__48817));
    LocalMux I__11004 (
            .O(N__48823),
            .I(N__48814));
    LocalMux I__11003 (
            .O(N__48820),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__11002 (
            .O(N__48817),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__11001 (
            .O(N__48814),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__11000 (
            .O(N__48807),
            .I(N__48804));
    LocalMux I__10999 (
            .O(N__48804),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__10998 (
            .O(N__48801),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__10997 (
            .O(N__48798),
            .I(N__48794));
    CascadeMux I__10996 (
            .O(N__48797),
            .I(N__48791));
    InMux I__10995 (
            .O(N__48794),
            .I(N__48788));
    InMux I__10994 (
            .O(N__48791),
            .I(N__48785));
    LocalMux I__10993 (
            .O(N__48788),
            .I(N__48779));
    LocalMux I__10992 (
            .O(N__48785),
            .I(N__48779));
    InMux I__10991 (
            .O(N__48784),
            .I(N__48776));
    Span4Mux_v I__10990 (
            .O(N__48779),
            .I(N__48773));
    LocalMux I__10989 (
            .O(N__48776),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__10988 (
            .O(N__48773),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__10987 (
            .O(N__48768),
            .I(bfn_17_22_0_));
    CascadeMux I__10986 (
            .O(N__48765),
            .I(N__48761));
    InMux I__10985 (
            .O(N__48764),
            .I(N__48758));
    InMux I__10984 (
            .O(N__48761),
            .I(N__48755));
    LocalMux I__10983 (
            .O(N__48758),
            .I(N__48751));
    LocalMux I__10982 (
            .O(N__48755),
            .I(N__48748));
    InMux I__10981 (
            .O(N__48754),
            .I(N__48745));
    Span4Mux_v I__10980 (
            .O(N__48751),
            .I(N__48740));
    Span4Mux_v I__10979 (
            .O(N__48748),
            .I(N__48740));
    LocalMux I__10978 (
            .O(N__48745),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__10977 (
            .O(N__48740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__10976 (
            .O(N__48735),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__10975 (
            .O(N__48732),
            .I(N__48729));
    InMux I__10974 (
            .O(N__48729),
            .I(N__48725));
    InMux I__10973 (
            .O(N__48728),
            .I(N__48722));
    LocalMux I__10972 (
            .O(N__48725),
            .I(N__48716));
    LocalMux I__10971 (
            .O(N__48722),
            .I(N__48716));
    InMux I__10970 (
            .O(N__48721),
            .I(N__48713));
    Span4Mux_h I__10969 (
            .O(N__48716),
            .I(N__48710));
    LocalMux I__10968 (
            .O(N__48713),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__10967 (
            .O(N__48710),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__10966 (
            .O(N__48705),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__10965 (
            .O(N__48702),
            .I(N__48698));
    CascadeMux I__10964 (
            .O(N__48701),
            .I(N__48695));
    InMux I__10963 (
            .O(N__48698),
            .I(N__48689));
    InMux I__10962 (
            .O(N__48695),
            .I(N__48689));
    InMux I__10961 (
            .O(N__48694),
            .I(N__48686));
    LocalMux I__10960 (
            .O(N__48689),
            .I(N__48683));
    LocalMux I__10959 (
            .O(N__48686),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv12 I__10958 (
            .O(N__48683),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__10957 (
            .O(N__48678),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__10956 (
            .O(N__48675),
            .I(N__48668));
    InMux I__10955 (
            .O(N__48674),
            .I(N__48668));
    InMux I__10954 (
            .O(N__48673),
            .I(N__48665));
    LocalMux I__10953 (
            .O(N__48668),
            .I(N__48662));
    LocalMux I__10952 (
            .O(N__48665),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv12 I__10951 (
            .O(N__48662),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__10950 (
            .O(N__48657),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__10949 (
            .O(N__48654),
            .I(N__48651));
    InMux I__10948 (
            .O(N__48651),
            .I(N__48646));
    InMux I__10947 (
            .O(N__48650),
            .I(N__48643));
    InMux I__10946 (
            .O(N__48649),
            .I(N__48640));
    LocalMux I__10945 (
            .O(N__48646),
            .I(N__48635));
    LocalMux I__10944 (
            .O(N__48643),
            .I(N__48635));
    LocalMux I__10943 (
            .O(N__48640),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv12 I__10942 (
            .O(N__48635),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__10941 (
            .O(N__48630),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__10940 (
            .O(N__48627),
            .I(N__48623));
    CascadeMux I__10939 (
            .O(N__48626),
            .I(N__48620));
    InMux I__10938 (
            .O(N__48623),
            .I(N__48614));
    InMux I__10937 (
            .O(N__48620),
            .I(N__48614));
    InMux I__10936 (
            .O(N__48619),
            .I(N__48611));
    LocalMux I__10935 (
            .O(N__48614),
            .I(N__48608));
    LocalMux I__10934 (
            .O(N__48611),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv12 I__10933 (
            .O(N__48608),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__10932 (
            .O(N__48603),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__10931 (
            .O(N__48600),
            .I(N__48593));
    InMux I__10930 (
            .O(N__48599),
            .I(N__48593));
    InMux I__10929 (
            .O(N__48598),
            .I(N__48590));
    LocalMux I__10928 (
            .O(N__48593),
            .I(N__48587));
    LocalMux I__10927 (
            .O(N__48590),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv12 I__10926 (
            .O(N__48587),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__10925 (
            .O(N__48582),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__10924 (
            .O(N__48579),
            .I(N__48575));
    CascadeMux I__10923 (
            .O(N__48578),
            .I(N__48572));
    InMux I__10922 (
            .O(N__48575),
            .I(N__48567));
    InMux I__10921 (
            .O(N__48572),
            .I(N__48567));
    LocalMux I__10920 (
            .O(N__48567),
            .I(N__48563));
    InMux I__10919 (
            .O(N__48566),
            .I(N__48560));
    Span4Mux_v I__10918 (
            .O(N__48563),
            .I(N__48557));
    LocalMux I__10917 (
            .O(N__48560),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__10916 (
            .O(N__48557),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__10915 (
            .O(N__48552),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__10914 (
            .O(N__48549),
            .I(N__48546));
    InMux I__10913 (
            .O(N__48546),
            .I(N__48543));
    LocalMux I__10912 (
            .O(N__48543),
            .I(N__48538));
    InMux I__10911 (
            .O(N__48542),
            .I(N__48535));
    InMux I__10910 (
            .O(N__48541),
            .I(N__48532));
    Span4Mux_h I__10909 (
            .O(N__48538),
            .I(N__48529));
    LocalMux I__10908 (
            .O(N__48535),
            .I(N__48526));
    LocalMux I__10907 (
            .O(N__48532),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__10906 (
            .O(N__48529),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv12 I__10905 (
            .O(N__48526),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__10904 (
            .O(N__48519),
            .I(bfn_17_21_0_));
    CascadeMux I__10903 (
            .O(N__48516),
            .I(N__48513));
    InMux I__10902 (
            .O(N__48513),
            .I(N__48509));
    InMux I__10901 (
            .O(N__48512),
            .I(N__48506));
    LocalMux I__10900 (
            .O(N__48509),
            .I(N__48500));
    LocalMux I__10899 (
            .O(N__48506),
            .I(N__48500));
    InMux I__10898 (
            .O(N__48505),
            .I(N__48497));
    Span4Mux_v I__10897 (
            .O(N__48500),
            .I(N__48494));
    LocalMux I__10896 (
            .O(N__48497),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__10895 (
            .O(N__48494),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__10894 (
            .O(N__48489),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__10893 (
            .O(N__48486),
            .I(N__48480));
    InMux I__10892 (
            .O(N__48485),
            .I(N__48480));
    LocalMux I__10891 (
            .O(N__48480),
            .I(N__48476));
    InMux I__10890 (
            .O(N__48479),
            .I(N__48473));
    Span4Mux_h I__10889 (
            .O(N__48476),
            .I(N__48470));
    LocalMux I__10888 (
            .O(N__48473),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__10887 (
            .O(N__48470),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__10886 (
            .O(N__48465),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__10885 (
            .O(N__48462),
            .I(N__48456));
    InMux I__10884 (
            .O(N__48461),
            .I(N__48456));
    LocalMux I__10883 (
            .O(N__48456),
            .I(N__48452));
    InMux I__10882 (
            .O(N__48455),
            .I(N__48449));
    Span4Mux_h I__10881 (
            .O(N__48452),
            .I(N__48446));
    LocalMux I__10880 (
            .O(N__48449),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__10879 (
            .O(N__48446),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__10878 (
            .O(N__48441),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__10877 (
            .O(N__48438),
            .I(N__48434));
    CascadeMux I__10876 (
            .O(N__48437),
            .I(N__48431));
    InMux I__10875 (
            .O(N__48434),
            .I(N__48426));
    InMux I__10874 (
            .O(N__48431),
            .I(N__48426));
    LocalMux I__10873 (
            .O(N__48426),
            .I(N__48422));
    InMux I__10872 (
            .O(N__48425),
            .I(N__48419));
    Span4Mux_v I__10871 (
            .O(N__48422),
            .I(N__48416));
    LocalMux I__10870 (
            .O(N__48419),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__10869 (
            .O(N__48416),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__10868 (
            .O(N__48411),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__10867 (
            .O(N__48408),
            .I(N__48404));
    CascadeMux I__10866 (
            .O(N__48407),
            .I(N__48401));
    InMux I__10865 (
            .O(N__48404),
            .I(N__48396));
    InMux I__10864 (
            .O(N__48401),
            .I(N__48396));
    LocalMux I__10863 (
            .O(N__48396),
            .I(N__48392));
    InMux I__10862 (
            .O(N__48395),
            .I(N__48389));
    Span4Mux_h I__10861 (
            .O(N__48392),
            .I(N__48386));
    LocalMux I__10860 (
            .O(N__48389),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__10859 (
            .O(N__48386),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__10858 (
            .O(N__48381),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__10857 (
            .O(N__48378),
            .I(N__48372));
    InMux I__10856 (
            .O(N__48377),
            .I(N__48372));
    LocalMux I__10855 (
            .O(N__48372),
            .I(N__48368));
    InMux I__10854 (
            .O(N__48371),
            .I(N__48365));
    Span4Mux_v I__10853 (
            .O(N__48368),
            .I(N__48362));
    LocalMux I__10852 (
            .O(N__48365),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__10851 (
            .O(N__48362),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__10850 (
            .O(N__48357),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__10849 (
            .O(N__48354),
            .I(N__48348));
    InMux I__10848 (
            .O(N__48353),
            .I(N__48348));
    LocalMux I__10847 (
            .O(N__48348),
            .I(N__48344));
    InMux I__10846 (
            .O(N__48347),
            .I(N__48341));
    Span4Mux_v I__10845 (
            .O(N__48344),
            .I(N__48338));
    LocalMux I__10844 (
            .O(N__48341),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__10843 (
            .O(N__48338),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__10842 (
            .O(N__48333),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__10841 (
            .O(N__48330),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__10840 (
            .O(N__48327),
            .I(N__48323));
    InMux I__10839 (
            .O(N__48326),
            .I(N__48320));
    LocalMux I__10838 (
            .O(N__48323),
            .I(N__48317));
    LocalMux I__10837 (
            .O(N__48320),
            .I(N__48314));
    Span4Mux_h I__10836 (
            .O(N__48317),
            .I(N__48309));
    Span4Mux_h I__10835 (
            .O(N__48314),
            .I(N__48309));
    Odrv4 I__10834 (
            .O(N__48309),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__10833 (
            .O(N__48306),
            .I(bfn_17_20_0_));
    InMux I__10832 (
            .O(N__48303),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__10831 (
            .O(N__48300),
            .I(N__48293));
    InMux I__10830 (
            .O(N__48299),
            .I(N__48293));
    InMux I__10829 (
            .O(N__48298),
            .I(N__48290));
    LocalMux I__10828 (
            .O(N__48293),
            .I(N__48287));
    LocalMux I__10827 (
            .O(N__48290),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv12 I__10826 (
            .O(N__48287),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__10825 (
            .O(N__48282),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__10824 (
            .O(N__48279),
            .I(N__48272));
    InMux I__10823 (
            .O(N__48278),
            .I(N__48272));
    InMux I__10822 (
            .O(N__48277),
            .I(N__48269));
    LocalMux I__10821 (
            .O(N__48272),
            .I(N__48266));
    LocalMux I__10820 (
            .O(N__48269),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv12 I__10819 (
            .O(N__48266),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__10818 (
            .O(N__48261),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__10817 (
            .O(N__48258),
            .I(N__48254));
    InMux I__10816 (
            .O(N__48257),
            .I(N__48250));
    InMux I__10815 (
            .O(N__48254),
            .I(N__48247));
    InMux I__10814 (
            .O(N__48253),
            .I(N__48244));
    LocalMux I__10813 (
            .O(N__48250),
            .I(N__48239));
    LocalMux I__10812 (
            .O(N__48247),
            .I(N__48239));
    LocalMux I__10811 (
            .O(N__48244),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv12 I__10810 (
            .O(N__48239),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__10809 (
            .O(N__48234),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__10808 (
            .O(N__48231),
            .I(N__48227));
    InMux I__10807 (
            .O(N__48230),
            .I(N__48224));
    InMux I__10806 (
            .O(N__48227),
            .I(N__48221));
    LocalMux I__10805 (
            .O(N__48224),
            .I(N__48217));
    LocalMux I__10804 (
            .O(N__48221),
            .I(N__48214));
    InMux I__10803 (
            .O(N__48220),
            .I(N__48211));
    Span4Mux_h I__10802 (
            .O(N__48217),
            .I(N__48206));
    Span4Mux_h I__10801 (
            .O(N__48214),
            .I(N__48206));
    LocalMux I__10800 (
            .O(N__48211),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__10799 (
            .O(N__48206),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__10798 (
            .O(N__48201),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__10797 (
            .O(N__48198),
            .I(N__48194));
    CascadeMux I__10796 (
            .O(N__48197),
            .I(N__48191));
    InMux I__10795 (
            .O(N__48194),
            .I(N__48186));
    InMux I__10794 (
            .O(N__48191),
            .I(N__48186));
    LocalMux I__10793 (
            .O(N__48186),
            .I(N__48182));
    InMux I__10792 (
            .O(N__48185),
            .I(N__48179));
    Span4Mux_v I__10791 (
            .O(N__48182),
            .I(N__48176));
    LocalMux I__10790 (
            .O(N__48179),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__10789 (
            .O(N__48176),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__10788 (
            .O(N__48171),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__10787 (
            .O(N__48168),
            .I(N__48164));
    CascadeMux I__10786 (
            .O(N__48167),
            .I(N__48161));
    LocalMux I__10785 (
            .O(N__48164),
            .I(N__48158));
    InMux I__10784 (
            .O(N__48161),
            .I(N__48155));
    Odrv4 I__10783 (
            .O(N__48158),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__10782 (
            .O(N__48155),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__10781 (
            .O(N__48150),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__10780 (
            .O(N__48147),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__10779 (
            .O(N__48144),
            .I(N__48141));
    LocalMux I__10778 (
            .O(N__48141),
            .I(N__48138));
    Span4Mux_h I__10777 (
            .O(N__48138),
            .I(N__48134));
    InMux I__10776 (
            .O(N__48137),
            .I(N__48131));
    Odrv4 I__10775 (
            .O(N__48134),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__10774 (
            .O(N__48131),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__10773 (
            .O(N__48126),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__10772 (
            .O(N__48123),
            .I(N__48119));
    InMux I__10771 (
            .O(N__48122),
            .I(N__48114));
    InMux I__10770 (
            .O(N__48119),
            .I(N__48114));
    LocalMux I__10769 (
            .O(N__48114),
            .I(N__48111));
    Odrv4 I__10768 (
            .O(N__48111),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__10767 (
            .O(N__48108),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__10766 (
            .O(N__48105),
            .I(N__48099));
    InMux I__10765 (
            .O(N__48104),
            .I(N__48099));
    LocalMux I__10764 (
            .O(N__48099),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__10763 (
            .O(N__48096),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__10762 (
            .O(N__48093),
            .I(bfn_17_19_0_));
    InMux I__10761 (
            .O(N__48090),
            .I(N__48087));
    LocalMux I__10760 (
            .O(N__48087),
            .I(N__48084));
    Span4Mux_v I__10759 (
            .O(N__48084),
            .I(N__48081));
    Span4Mux_v I__10758 (
            .O(N__48081),
            .I(N__48077));
    InMux I__10757 (
            .O(N__48080),
            .I(N__48074));
    Odrv4 I__10756 (
            .O(N__48077),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__10755 (
            .O(N__48074),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__10754 (
            .O(N__48069),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__10753 (
            .O(N__48066),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__10752 (
            .O(N__48063),
            .I(N__48060));
    LocalMux I__10751 (
            .O(N__48060),
            .I(N__48056));
    CascadeMux I__10750 (
            .O(N__48059),
            .I(N__48053));
    Span4Mux_h I__10749 (
            .O(N__48056),
            .I(N__48050));
    InMux I__10748 (
            .O(N__48053),
            .I(N__48047));
    Odrv4 I__10747 (
            .O(N__48050),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__10746 (
            .O(N__48047),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__10745 (
            .O(N__48042),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__10744 (
            .O(N__48039),
            .I(N__48036));
    LocalMux I__10743 (
            .O(N__48036),
            .I(N__48033));
    Span4Mux_h I__10742 (
            .O(N__48033),
            .I(N__48029));
    InMux I__10741 (
            .O(N__48032),
            .I(N__48026));
    Odrv4 I__10740 (
            .O(N__48029),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__10739 (
            .O(N__48026),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__10738 (
            .O(N__48021),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__10737 (
            .O(N__48018),
            .I(N__48015));
    LocalMux I__10736 (
            .O(N__48015),
            .I(N__48011));
    InMux I__10735 (
            .O(N__48014),
            .I(N__48008));
    Odrv4 I__10734 (
            .O(N__48011),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__10733 (
            .O(N__48008),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__10732 (
            .O(N__48003),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__10731 (
            .O(N__48000),
            .I(N__47997));
    LocalMux I__10730 (
            .O(N__47997),
            .I(N__47994));
    Span4Mux_h I__10729 (
            .O(N__47994),
            .I(N__47990));
    InMux I__10728 (
            .O(N__47993),
            .I(N__47987));
    Odrv4 I__10727 (
            .O(N__47990),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__10726 (
            .O(N__47987),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__10725 (
            .O(N__47982),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__10724 (
            .O(N__47979),
            .I(N__47976));
    LocalMux I__10723 (
            .O(N__47976),
            .I(N__47972));
    InMux I__10722 (
            .O(N__47975),
            .I(N__47969));
    Odrv4 I__10721 (
            .O(N__47972),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__10720 (
            .O(N__47969),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__10719 (
            .O(N__47964),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__10718 (
            .O(N__47961),
            .I(N__47958));
    LocalMux I__10717 (
            .O(N__47958),
            .I(N__47954));
    CascadeMux I__10716 (
            .O(N__47957),
            .I(N__47951));
    Span4Mux_v I__10715 (
            .O(N__47954),
            .I(N__47948));
    InMux I__10714 (
            .O(N__47951),
            .I(N__47945));
    Odrv4 I__10713 (
            .O(N__47948),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__10712 (
            .O(N__47945),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__10711 (
            .O(N__47940),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__10710 (
            .O(N__47937),
            .I(N__47934));
    LocalMux I__10709 (
            .O(N__47934),
            .I(N__47931));
    Span4Mux_h I__10708 (
            .O(N__47931),
            .I(N__47927));
    InMux I__10707 (
            .O(N__47930),
            .I(N__47924));
    Odrv4 I__10706 (
            .O(N__47927),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    LocalMux I__10705 (
            .O(N__47924),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__10704 (
            .O(N__47919),
            .I(bfn_17_18_0_));
    InMux I__10703 (
            .O(N__47916),
            .I(N__47913));
    LocalMux I__10702 (
            .O(N__47913),
            .I(N__47910));
    Span4Mux_h I__10701 (
            .O(N__47910),
            .I(N__47906));
    InMux I__10700 (
            .O(N__47909),
            .I(N__47903));
    Odrv4 I__10699 (
            .O(N__47906),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__10698 (
            .O(N__47903),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__10697 (
            .O(N__47898),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__10696 (
            .O(N__47895),
            .I(N__47891));
    InMux I__10695 (
            .O(N__47894),
            .I(N__47888));
    LocalMux I__10694 (
            .O(N__47891),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__10693 (
            .O(N__47888),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__10692 (
            .O(N__47883),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__10691 (
            .O(N__47880),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__10690 (
            .O(N__47877),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__10689 (
            .O(N__47874),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__10688 (
            .O(N__47871),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__10687 (
            .O(N__47868),
            .I(N__47865));
    LocalMux I__10686 (
            .O(N__47865),
            .I(N__47862));
    Span4Mux_h I__10685 (
            .O(N__47862),
            .I(N__47858));
    InMux I__10684 (
            .O(N__47861),
            .I(N__47855));
    Odrv4 I__10683 (
            .O(N__47858),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    LocalMux I__10682 (
            .O(N__47855),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__10681 (
            .O(N__47850),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__10680 (
            .O(N__47847),
            .I(N__47844));
    LocalMux I__10679 (
            .O(N__47844),
            .I(N__47841));
    Span4Mux_h I__10678 (
            .O(N__47841),
            .I(N__47837));
    InMux I__10677 (
            .O(N__47840),
            .I(N__47834));
    Odrv4 I__10676 (
            .O(N__47837),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__10675 (
            .O(N__47834),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__10674 (
            .O(N__47829),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__10673 (
            .O(N__47826),
            .I(N__47823));
    LocalMux I__10672 (
            .O(N__47823),
            .I(N__47819));
    InMux I__10671 (
            .O(N__47822),
            .I(N__47816));
    Odrv4 I__10670 (
            .O(N__47819),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__10669 (
            .O(N__47816),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__10668 (
            .O(N__47811),
            .I(bfn_17_17_0_));
    InMux I__10667 (
            .O(N__47808),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__10666 (
            .O(N__47805),
            .I(N__47802));
    LocalMux I__10665 (
            .O(N__47802),
            .I(N__47799));
    Odrv4 I__10664 (
            .O(N__47799),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ));
    InMux I__10663 (
            .O(N__47796),
            .I(N__47792));
    InMux I__10662 (
            .O(N__47795),
            .I(N__47789));
    LocalMux I__10661 (
            .O(N__47792),
            .I(N__47784));
    LocalMux I__10660 (
            .O(N__47789),
            .I(N__47784));
    Span4Mux_v I__10659 (
            .O(N__47784),
            .I(N__47781));
    Odrv4 I__10658 (
            .O(N__47781),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ));
    InMux I__10657 (
            .O(N__47778),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ));
    InMux I__10656 (
            .O(N__47775),
            .I(N__47771));
    InMux I__10655 (
            .O(N__47774),
            .I(N__47768));
    LocalMux I__10654 (
            .O(N__47771),
            .I(N__47763));
    LocalMux I__10653 (
            .O(N__47768),
            .I(N__47763));
    Odrv12 I__10652 (
            .O(N__47763),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ));
    InMux I__10651 (
            .O(N__47760),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ));
    InMux I__10650 (
            .O(N__47757),
            .I(N__47754));
    LocalMux I__10649 (
            .O(N__47754),
            .I(N__47751));
    Span4Mux_v I__10648 (
            .O(N__47751),
            .I(N__47748));
    Odrv4 I__10647 (
            .O(N__47748),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ));
    InMux I__10646 (
            .O(N__47745),
            .I(N__47741));
    InMux I__10645 (
            .O(N__47744),
            .I(N__47738));
    LocalMux I__10644 (
            .O(N__47741),
            .I(N__47733));
    LocalMux I__10643 (
            .O(N__47738),
            .I(N__47733));
    Odrv12 I__10642 (
            .O(N__47733),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ));
    InMux I__10641 (
            .O(N__47730),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ));
    InMux I__10640 (
            .O(N__47727),
            .I(N__47723));
    InMux I__10639 (
            .O(N__47726),
            .I(N__47720));
    LocalMux I__10638 (
            .O(N__47723),
            .I(N__47715));
    LocalMux I__10637 (
            .O(N__47720),
            .I(N__47715));
    Span4Mux_v I__10636 (
            .O(N__47715),
            .I(N__47712));
    Odrv4 I__10635 (
            .O(N__47712),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ));
    InMux I__10634 (
            .O(N__47709),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ));
    InMux I__10633 (
            .O(N__47706),
            .I(N__47703));
    LocalMux I__10632 (
            .O(N__47703),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ));
    InMux I__10631 (
            .O(N__47700),
            .I(N__47696));
    InMux I__10630 (
            .O(N__47699),
            .I(N__47693));
    LocalMux I__10629 (
            .O(N__47696),
            .I(N__47688));
    LocalMux I__10628 (
            .O(N__47693),
            .I(N__47688));
    Odrv12 I__10627 (
            .O(N__47688),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ));
    InMux I__10626 (
            .O(N__47685),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ));
    InMux I__10625 (
            .O(N__47682),
            .I(N__47679));
    LocalMux I__10624 (
            .O(N__47679),
            .I(N__47676));
    Span4Mux_v I__10623 (
            .O(N__47676),
            .I(N__47673));
    Odrv4 I__10622 (
            .O(N__47673),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ));
    InMux I__10621 (
            .O(N__47670),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ));
    InMux I__10620 (
            .O(N__47667),
            .I(N__47664));
    LocalMux I__10619 (
            .O(N__47664),
            .I(N__47661));
    Span4Mux_h I__10618 (
            .O(N__47661),
            .I(N__47657));
    InMux I__10617 (
            .O(N__47660),
            .I(N__47654));
    Span4Mux_v I__10616 (
            .O(N__47657),
            .I(N__47651));
    LocalMux I__10615 (
            .O(N__47654),
            .I(N__47648));
    Odrv4 I__10614 (
            .O(N__47651),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_28));
    Odrv12 I__10613 (
            .O(N__47648),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_28));
    InMux I__10612 (
            .O(N__47643),
            .I(N__47639));
    InMux I__10611 (
            .O(N__47642),
            .I(N__47636));
    LocalMux I__10610 (
            .O(N__47639),
            .I(N__47632));
    LocalMux I__10609 (
            .O(N__47636),
            .I(N__47629));
    InMux I__10608 (
            .O(N__47635),
            .I(N__47626));
    Span4Mux_h I__10607 (
            .O(N__47632),
            .I(N__47622));
    Span4Mux_h I__10606 (
            .O(N__47629),
            .I(N__47619));
    LocalMux I__10605 (
            .O(N__47626),
            .I(N__47614));
    InMux I__10604 (
            .O(N__47625),
            .I(N__47611));
    Span4Mux_v I__10603 (
            .O(N__47622),
            .I(N__47608));
    Span4Mux_h I__10602 (
            .O(N__47619),
            .I(N__47605));
    InMux I__10601 (
            .O(N__47618),
            .I(N__47600));
    InMux I__10600 (
            .O(N__47617),
            .I(N__47600));
    Span12Mux_s9_v I__10599 (
            .O(N__47614),
            .I(N__47595));
    LocalMux I__10598 (
            .O(N__47611),
            .I(N__47595));
    Odrv4 I__10597 (
            .O(N__47608),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__10596 (
            .O(N__47605),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__10595 (
            .O(N__47600),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv12 I__10594 (
            .O(N__47595),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__10593 (
            .O(N__47586),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__10592 (
            .O(N__47583),
            .I(N__47580));
    LocalMux I__10591 (
            .O(N__47580),
            .I(N__47577));
    Odrv4 I__10590 (
            .O(N__47577),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ));
    InMux I__10589 (
            .O(N__47574),
            .I(N__47570));
    InMux I__10588 (
            .O(N__47573),
            .I(N__47567));
    LocalMux I__10587 (
            .O(N__47570),
            .I(N__47562));
    LocalMux I__10586 (
            .O(N__47567),
            .I(N__47562));
    Span4Mux_v I__10585 (
            .O(N__47562),
            .I(N__47559));
    Odrv4 I__10584 (
            .O(N__47559),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ));
    InMux I__10583 (
            .O(N__47556),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ));
    InMux I__10582 (
            .O(N__47553),
            .I(N__47550));
    LocalMux I__10581 (
            .O(N__47550),
            .I(N__47547));
    Span4Mux_h I__10580 (
            .O(N__47547),
            .I(N__47544));
    Odrv4 I__10579 (
            .O(N__47544),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ));
    InMux I__10578 (
            .O(N__47541),
            .I(N__47537));
    InMux I__10577 (
            .O(N__47540),
            .I(N__47534));
    LocalMux I__10576 (
            .O(N__47537),
            .I(N__47529));
    LocalMux I__10575 (
            .O(N__47534),
            .I(N__47529));
    Span4Mux_h I__10574 (
            .O(N__47529),
            .I(N__47526));
    Odrv4 I__10573 (
            .O(N__47526),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ));
    InMux I__10572 (
            .O(N__47523),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ));
    InMux I__10571 (
            .O(N__47520),
            .I(N__47517));
    LocalMux I__10570 (
            .O(N__47517),
            .I(N__47514));
    Odrv4 I__10569 (
            .O(N__47514),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ));
    InMux I__10568 (
            .O(N__47511),
            .I(N__47507));
    InMux I__10567 (
            .O(N__47510),
            .I(N__47504));
    LocalMux I__10566 (
            .O(N__47507),
            .I(N__47499));
    LocalMux I__10565 (
            .O(N__47504),
            .I(N__47499));
    Span4Mux_h I__10564 (
            .O(N__47499),
            .I(N__47496));
    Odrv4 I__10563 (
            .O(N__47496),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ));
    InMux I__10562 (
            .O(N__47493),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ));
    InMux I__10561 (
            .O(N__47490),
            .I(N__47487));
    LocalMux I__10560 (
            .O(N__47487),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ));
    InMux I__10559 (
            .O(N__47484),
            .I(N__47480));
    InMux I__10558 (
            .O(N__47483),
            .I(N__47477));
    LocalMux I__10557 (
            .O(N__47480),
            .I(N__47472));
    LocalMux I__10556 (
            .O(N__47477),
            .I(N__47472));
    Odrv12 I__10555 (
            .O(N__47472),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ));
    InMux I__10554 (
            .O(N__47469),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ));
    InMux I__10553 (
            .O(N__47466),
            .I(N__47463));
    LocalMux I__10552 (
            .O(N__47463),
            .I(N__47460));
    Odrv4 I__10551 (
            .O(N__47460),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ));
    InMux I__10550 (
            .O(N__47457),
            .I(N__47453));
    InMux I__10549 (
            .O(N__47456),
            .I(N__47450));
    LocalMux I__10548 (
            .O(N__47453),
            .I(N__47445));
    LocalMux I__10547 (
            .O(N__47450),
            .I(N__47445));
    Span4Mux_h I__10546 (
            .O(N__47445),
            .I(N__47442));
    Odrv4 I__10545 (
            .O(N__47442),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ));
    InMux I__10544 (
            .O(N__47439),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ));
    InMux I__10543 (
            .O(N__47436),
            .I(N__47432));
    InMux I__10542 (
            .O(N__47435),
            .I(N__47429));
    LocalMux I__10541 (
            .O(N__47432),
            .I(N__47424));
    LocalMux I__10540 (
            .O(N__47429),
            .I(N__47424));
    Odrv12 I__10539 (
            .O(N__47424),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ));
    InMux I__10538 (
            .O(N__47421),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ));
    InMux I__10537 (
            .O(N__47418),
            .I(N__47415));
    LocalMux I__10536 (
            .O(N__47415),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ));
    InMux I__10535 (
            .O(N__47412),
            .I(N__47408));
    InMux I__10534 (
            .O(N__47411),
            .I(N__47405));
    LocalMux I__10533 (
            .O(N__47408),
            .I(N__47400));
    LocalMux I__10532 (
            .O(N__47405),
            .I(N__47400));
    Odrv12 I__10531 (
            .O(N__47400),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ));
    InMux I__10530 (
            .O(N__47397),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ));
    InMux I__10529 (
            .O(N__47394),
            .I(N__47391));
    LocalMux I__10528 (
            .O(N__47391),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ));
    InMux I__10527 (
            .O(N__47388),
            .I(N__47384));
    InMux I__10526 (
            .O(N__47387),
            .I(N__47381));
    LocalMux I__10525 (
            .O(N__47384),
            .I(N__47376));
    LocalMux I__10524 (
            .O(N__47381),
            .I(N__47376));
    Span4Mux_v I__10523 (
            .O(N__47376),
            .I(N__47373));
    Odrv4 I__10522 (
            .O(N__47373),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ));
    InMux I__10521 (
            .O(N__47370),
            .I(bfn_17_15_0_));
    InMux I__10520 (
            .O(N__47367),
            .I(N__47364));
    LocalMux I__10519 (
            .O(N__47364),
            .I(N__47360));
    InMux I__10518 (
            .O(N__47363),
            .I(N__47357));
    Span4Mux_v I__10517 (
            .O(N__47360),
            .I(N__47354));
    LocalMux I__10516 (
            .O(N__47357),
            .I(N__47351));
    Odrv4 I__10515 (
            .O(N__47354),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ));
    Odrv12 I__10514 (
            .O(N__47351),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ));
    InMux I__10513 (
            .O(N__47346),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ));
    InMux I__10512 (
            .O(N__47343),
            .I(N__47340));
    LocalMux I__10511 (
            .O(N__47340),
            .I(N__47337));
    Odrv4 I__10510 (
            .O(N__47337),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ));
    InMux I__10509 (
            .O(N__47334),
            .I(N__47330));
    InMux I__10508 (
            .O(N__47333),
            .I(N__47327));
    LocalMux I__10507 (
            .O(N__47330),
            .I(N__47322));
    LocalMux I__10506 (
            .O(N__47327),
            .I(N__47322));
    Span4Mux_h I__10505 (
            .O(N__47322),
            .I(N__47319));
    Odrv4 I__10504 (
            .O(N__47319),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ));
    InMux I__10503 (
            .O(N__47316),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ));
    InMux I__10502 (
            .O(N__47313),
            .I(N__47309));
    InMux I__10501 (
            .O(N__47312),
            .I(N__47306));
    LocalMux I__10500 (
            .O(N__47309),
            .I(N__47301));
    LocalMux I__10499 (
            .O(N__47306),
            .I(N__47301));
    Span4Mux_h I__10498 (
            .O(N__47301),
            .I(N__47298));
    Odrv4 I__10497 (
            .O(N__47298),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ));
    InMux I__10496 (
            .O(N__47295),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ));
    InMux I__10495 (
            .O(N__47292),
            .I(N__47288));
    InMux I__10494 (
            .O(N__47291),
            .I(N__47285));
    LocalMux I__10493 (
            .O(N__47288),
            .I(N__47282));
    LocalMux I__10492 (
            .O(N__47285),
            .I(N__47279));
    Span4Mux_v I__10491 (
            .O(N__47282),
            .I(N__47274));
    Span4Mux_v I__10490 (
            .O(N__47279),
            .I(N__47274));
    Odrv4 I__10489 (
            .O(N__47274),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ));
    InMux I__10488 (
            .O(N__47271),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ));
    InMux I__10487 (
            .O(N__47268),
            .I(N__47265));
    LocalMux I__10486 (
            .O(N__47265),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ));
    InMux I__10485 (
            .O(N__47262),
            .I(N__47258));
    InMux I__10484 (
            .O(N__47261),
            .I(N__47255));
    LocalMux I__10483 (
            .O(N__47258),
            .I(N__47250));
    LocalMux I__10482 (
            .O(N__47255),
            .I(N__47250));
    Span4Mux_h I__10481 (
            .O(N__47250),
            .I(N__47247));
    Odrv4 I__10480 (
            .O(N__47247),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ));
    InMux I__10479 (
            .O(N__47244),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ));
    InMux I__10478 (
            .O(N__47241),
            .I(N__47238));
    LocalMux I__10477 (
            .O(N__47238),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ));
    InMux I__10476 (
            .O(N__47235),
            .I(N__47231));
    InMux I__10475 (
            .O(N__47234),
            .I(N__47228));
    LocalMux I__10474 (
            .O(N__47231),
            .I(N__47223));
    LocalMux I__10473 (
            .O(N__47228),
            .I(N__47223));
    Odrv12 I__10472 (
            .O(N__47223),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ));
    InMux I__10471 (
            .O(N__47220),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ));
    InMux I__10470 (
            .O(N__47217),
            .I(N__47214));
    LocalMux I__10469 (
            .O(N__47214),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ));
    InMux I__10468 (
            .O(N__47211),
            .I(N__47207));
    InMux I__10467 (
            .O(N__47210),
            .I(N__47204));
    LocalMux I__10466 (
            .O(N__47207),
            .I(N__47199));
    LocalMux I__10465 (
            .O(N__47204),
            .I(N__47199));
    Span4Mux_h I__10464 (
            .O(N__47199),
            .I(N__47196));
    Span4Mux_v I__10463 (
            .O(N__47196),
            .I(N__47193));
    Odrv4 I__10462 (
            .O(N__47193),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ));
    InMux I__10461 (
            .O(N__47190),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ));
    InMux I__10460 (
            .O(N__47187),
            .I(N__47184));
    LocalMux I__10459 (
            .O(N__47184),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ));
    InMux I__10458 (
            .O(N__47181),
            .I(N__47177));
    InMux I__10457 (
            .O(N__47180),
            .I(N__47174));
    LocalMux I__10456 (
            .O(N__47177),
            .I(N__47169));
    LocalMux I__10455 (
            .O(N__47174),
            .I(N__47169));
    Odrv12 I__10454 (
            .O(N__47169),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ));
    InMux I__10453 (
            .O(N__47166),
            .I(bfn_17_14_0_));
    InMux I__10452 (
            .O(N__47163),
            .I(N__47160));
    LocalMux I__10451 (
            .O(N__47160),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ));
    InMux I__10450 (
            .O(N__47157),
            .I(N__47154));
    LocalMux I__10449 (
            .O(N__47154),
            .I(N__47150));
    CascadeMux I__10448 (
            .O(N__47153),
            .I(N__47146));
    Span4Mux_v I__10447 (
            .O(N__47150),
            .I(N__47143));
    InMux I__10446 (
            .O(N__47149),
            .I(N__47140));
    InMux I__10445 (
            .O(N__47146),
            .I(N__47137));
    Span4Mux_h I__10444 (
            .O(N__47143),
            .I(N__47134));
    LocalMux I__10443 (
            .O(N__47140),
            .I(N__47131));
    LocalMux I__10442 (
            .O(N__47137),
            .I(N__47128));
    Span4Mux_h I__10441 (
            .O(N__47134),
            .I(N__47125));
    Span4Mux_h I__10440 (
            .O(N__47131),
            .I(N__47120));
    Span4Mux_h I__10439 (
            .O(N__47128),
            .I(N__47120));
    Odrv4 I__10438 (
            .O(N__47125),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    Odrv4 I__10437 (
            .O(N__47120),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    InMux I__10436 (
            .O(N__47115),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ));
    InMux I__10435 (
            .O(N__47112),
            .I(N__47109));
    LocalMux I__10434 (
            .O(N__47109),
            .I(N__47106));
    Odrv4 I__10433 (
            .O(N__47106),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ));
    InMux I__10432 (
            .O(N__47103),
            .I(N__47099));
    InMux I__10431 (
            .O(N__47102),
            .I(N__47096));
    LocalMux I__10430 (
            .O(N__47099),
            .I(N__47091));
    LocalMux I__10429 (
            .O(N__47096),
            .I(N__47091));
    Span4Mux_v I__10428 (
            .O(N__47091),
            .I(N__47088));
    Odrv4 I__10427 (
            .O(N__47088),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ));
    InMux I__10426 (
            .O(N__47085),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ));
    InMux I__10425 (
            .O(N__47082),
            .I(N__47078));
    InMux I__10424 (
            .O(N__47081),
            .I(N__47075));
    LocalMux I__10423 (
            .O(N__47078),
            .I(N__47070));
    LocalMux I__10422 (
            .O(N__47075),
            .I(N__47070));
    Odrv12 I__10421 (
            .O(N__47070),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ));
    InMux I__10420 (
            .O(N__47067),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ));
    InMux I__10419 (
            .O(N__47064),
            .I(N__47061));
    LocalMux I__10418 (
            .O(N__47061),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ));
    InMux I__10417 (
            .O(N__47058),
            .I(N__47054));
    InMux I__10416 (
            .O(N__47057),
            .I(N__47051));
    LocalMux I__10415 (
            .O(N__47054),
            .I(N__47046));
    LocalMux I__10414 (
            .O(N__47051),
            .I(N__47046));
    Odrv12 I__10413 (
            .O(N__47046),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ));
    InMux I__10412 (
            .O(N__47043),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ));
    InMux I__10411 (
            .O(N__47040),
            .I(N__47037));
    LocalMux I__10410 (
            .O(N__47037),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ));
    InMux I__10409 (
            .O(N__47034),
            .I(N__47030));
    InMux I__10408 (
            .O(N__47033),
            .I(N__47027));
    LocalMux I__10407 (
            .O(N__47030),
            .I(N__47022));
    LocalMux I__10406 (
            .O(N__47027),
            .I(N__47022));
    Span4Mux_v I__10405 (
            .O(N__47022),
            .I(N__47019));
    Odrv4 I__10404 (
            .O(N__47019),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ));
    InMux I__10403 (
            .O(N__47016),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ));
    InMux I__10402 (
            .O(N__47013),
            .I(N__47010));
    LocalMux I__10401 (
            .O(N__47010),
            .I(N__47007));
    Span4Mux_h I__10400 (
            .O(N__47007),
            .I(N__47004));
    Odrv4 I__10399 (
            .O(N__47004),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ));
    InMux I__10398 (
            .O(N__47001),
            .I(N__46997));
    InMux I__10397 (
            .O(N__47000),
            .I(N__46994));
    LocalMux I__10396 (
            .O(N__46997),
            .I(N__46989));
    LocalMux I__10395 (
            .O(N__46994),
            .I(N__46989));
    Span4Mux_v I__10394 (
            .O(N__46989),
            .I(N__46986));
    Odrv4 I__10393 (
            .O(N__46986),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ));
    InMux I__10392 (
            .O(N__46983),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ));
    InMux I__10391 (
            .O(N__46980),
            .I(N__46977));
    LocalMux I__10390 (
            .O(N__46977),
            .I(N__46974));
    Span4Mux_v I__10389 (
            .O(N__46974),
            .I(N__46971));
    Odrv4 I__10388 (
            .O(N__46971),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ));
    InMux I__10387 (
            .O(N__46968),
            .I(N__46964));
    InMux I__10386 (
            .O(N__46967),
            .I(N__46961));
    LocalMux I__10385 (
            .O(N__46964),
            .I(N__46956));
    LocalMux I__10384 (
            .O(N__46961),
            .I(N__46956));
    Odrv12 I__10383 (
            .O(N__46956),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ));
    InMux I__10382 (
            .O(N__46953),
            .I(bfn_17_13_0_));
    InMux I__10381 (
            .O(N__46950),
            .I(N__46947));
    LocalMux I__10380 (
            .O(N__46947),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ));
    InMux I__10379 (
            .O(N__46944),
            .I(N__46941));
    LocalMux I__10378 (
            .O(N__46941),
            .I(N__46937));
    InMux I__10377 (
            .O(N__46940),
            .I(N__46934));
    Span4Mux_v I__10376 (
            .O(N__46937),
            .I(N__46929));
    LocalMux I__10375 (
            .O(N__46934),
            .I(N__46929));
    Odrv4 I__10374 (
            .O(N__46929),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_22));
    InMux I__10373 (
            .O(N__46926),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ));
    InMux I__10372 (
            .O(N__46923),
            .I(N__46919));
    InMux I__10371 (
            .O(N__46922),
            .I(N__46916));
    LocalMux I__10370 (
            .O(N__46919),
            .I(N__46913));
    LocalMux I__10369 (
            .O(N__46916),
            .I(N__46910));
    Span4Mux_h I__10368 (
            .O(N__46913),
            .I(N__46907));
    Span4Mux_h I__10367 (
            .O(N__46910),
            .I(N__46904));
    Odrv4 I__10366 (
            .O(N__46907),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_23));
    Odrv4 I__10365 (
            .O(N__46904),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_23));
    InMux I__10364 (
            .O(N__46899),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ));
    InMux I__10363 (
            .O(N__46896),
            .I(bfn_17_11_0_));
    InMux I__10362 (
            .O(N__46893),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ));
    InMux I__10361 (
            .O(N__46890),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ));
    CascadeMux I__10360 (
            .O(N__46887),
            .I(N__46869));
    CascadeMux I__10359 (
            .O(N__46886),
            .I(N__46866));
    CascadeMux I__10358 (
            .O(N__46885),
            .I(N__46863));
    CascadeMux I__10357 (
            .O(N__46884),
            .I(N__46860));
    CascadeMux I__10356 (
            .O(N__46883),
            .I(N__46857));
    CascadeMux I__10355 (
            .O(N__46882),
            .I(N__46854));
    CascadeMux I__10354 (
            .O(N__46881),
            .I(N__46833));
    CascadeMux I__10353 (
            .O(N__46880),
            .I(N__46830));
    CascadeMux I__10352 (
            .O(N__46879),
            .I(N__46825));
    CascadeMux I__10351 (
            .O(N__46878),
            .I(N__46822));
    CascadeMux I__10350 (
            .O(N__46877),
            .I(N__46819));
    CascadeMux I__10349 (
            .O(N__46876),
            .I(N__46816));
    CascadeMux I__10348 (
            .O(N__46875),
            .I(N__46813));
    CascadeMux I__10347 (
            .O(N__46874),
            .I(N__46810));
    CascadeMux I__10346 (
            .O(N__46873),
            .I(N__46807));
    CascadeMux I__10345 (
            .O(N__46872),
            .I(N__46804));
    InMux I__10344 (
            .O(N__46869),
            .I(N__46799));
    InMux I__10343 (
            .O(N__46866),
            .I(N__46799));
    InMux I__10342 (
            .O(N__46863),
            .I(N__46790));
    InMux I__10341 (
            .O(N__46860),
            .I(N__46790));
    InMux I__10340 (
            .O(N__46857),
            .I(N__46790));
    InMux I__10339 (
            .O(N__46854),
            .I(N__46790));
    CascadeMux I__10338 (
            .O(N__46853),
            .I(N__46787));
    CascadeMux I__10337 (
            .O(N__46852),
            .I(N__46784));
    CascadeMux I__10336 (
            .O(N__46851),
            .I(N__46781));
    CascadeMux I__10335 (
            .O(N__46850),
            .I(N__46778));
    CascadeMux I__10334 (
            .O(N__46849),
            .I(N__46775));
    CascadeMux I__10333 (
            .O(N__46848),
            .I(N__46772));
    CascadeMux I__10332 (
            .O(N__46847),
            .I(N__46754));
    CascadeMux I__10331 (
            .O(N__46846),
            .I(N__46751));
    CascadeMux I__10330 (
            .O(N__46845),
            .I(N__46748));
    CascadeMux I__10329 (
            .O(N__46844),
            .I(N__46745));
    CascadeMux I__10328 (
            .O(N__46843),
            .I(N__46742));
    CascadeMux I__10327 (
            .O(N__46842),
            .I(N__46739));
    CascadeMux I__10326 (
            .O(N__46841),
            .I(N__46736));
    CascadeMux I__10325 (
            .O(N__46840),
            .I(N__46733));
    CascadeMux I__10324 (
            .O(N__46839),
            .I(N__46730));
    CascadeMux I__10323 (
            .O(N__46838),
            .I(N__46727));
    CascadeMux I__10322 (
            .O(N__46837),
            .I(N__46724));
    CascadeMux I__10321 (
            .O(N__46836),
            .I(N__46721));
    InMux I__10320 (
            .O(N__46833),
            .I(N__46718));
    InMux I__10319 (
            .O(N__46830),
            .I(N__46713));
    InMux I__10318 (
            .O(N__46829),
            .I(N__46713));
    InMux I__10317 (
            .O(N__46828),
            .I(N__46710));
    InMux I__10316 (
            .O(N__46825),
            .I(N__46705));
    InMux I__10315 (
            .O(N__46822),
            .I(N__46705));
    InMux I__10314 (
            .O(N__46819),
            .I(N__46700));
    InMux I__10313 (
            .O(N__46816),
            .I(N__46700));
    InMux I__10312 (
            .O(N__46813),
            .I(N__46691));
    InMux I__10311 (
            .O(N__46810),
            .I(N__46691));
    InMux I__10310 (
            .O(N__46807),
            .I(N__46691));
    InMux I__10309 (
            .O(N__46804),
            .I(N__46691));
    LocalMux I__10308 (
            .O(N__46799),
            .I(N__46681));
    LocalMux I__10307 (
            .O(N__46790),
            .I(N__46678));
    InMux I__10306 (
            .O(N__46787),
            .I(N__46669));
    InMux I__10305 (
            .O(N__46784),
            .I(N__46669));
    InMux I__10304 (
            .O(N__46781),
            .I(N__46669));
    InMux I__10303 (
            .O(N__46778),
            .I(N__46669));
    InMux I__10302 (
            .O(N__46775),
            .I(N__46664));
    InMux I__10301 (
            .O(N__46772),
            .I(N__46664));
    CascadeMux I__10300 (
            .O(N__46771),
            .I(N__46661));
    CascadeMux I__10299 (
            .O(N__46770),
            .I(N__46658));
    CascadeMux I__10298 (
            .O(N__46769),
            .I(N__46655));
    CascadeMux I__10297 (
            .O(N__46768),
            .I(N__46652));
    CascadeMux I__10296 (
            .O(N__46767),
            .I(N__46649));
    CascadeMux I__10295 (
            .O(N__46766),
            .I(N__46646));
    CascadeMux I__10294 (
            .O(N__46765),
            .I(N__46643));
    CascadeMux I__10293 (
            .O(N__46764),
            .I(N__46640));
    CascadeMux I__10292 (
            .O(N__46763),
            .I(N__46637));
    CascadeMux I__10291 (
            .O(N__46762),
            .I(N__46634));
    CascadeMux I__10290 (
            .O(N__46761),
            .I(N__46631));
    CascadeMux I__10289 (
            .O(N__46760),
            .I(N__46628));
    CascadeMux I__10288 (
            .O(N__46759),
            .I(N__46625));
    CascadeMux I__10287 (
            .O(N__46758),
            .I(N__46622));
    CascadeMux I__10286 (
            .O(N__46757),
            .I(N__46619));
    InMux I__10285 (
            .O(N__46754),
            .I(N__46610));
    InMux I__10284 (
            .O(N__46751),
            .I(N__46610));
    InMux I__10283 (
            .O(N__46748),
            .I(N__46610));
    InMux I__10282 (
            .O(N__46745),
            .I(N__46610));
    InMux I__10281 (
            .O(N__46742),
            .I(N__46601));
    InMux I__10280 (
            .O(N__46739),
            .I(N__46601));
    InMux I__10279 (
            .O(N__46736),
            .I(N__46601));
    InMux I__10278 (
            .O(N__46733),
            .I(N__46601));
    InMux I__10277 (
            .O(N__46730),
            .I(N__46592));
    InMux I__10276 (
            .O(N__46727),
            .I(N__46592));
    InMux I__10275 (
            .O(N__46724),
            .I(N__46592));
    InMux I__10274 (
            .O(N__46721),
            .I(N__46592));
    LocalMux I__10273 (
            .O(N__46718),
            .I(N__46587));
    LocalMux I__10272 (
            .O(N__46713),
            .I(N__46587));
    LocalMux I__10271 (
            .O(N__46710),
            .I(N__46573));
    LocalMux I__10270 (
            .O(N__46705),
            .I(N__46566));
    LocalMux I__10269 (
            .O(N__46700),
            .I(N__46566));
    LocalMux I__10268 (
            .O(N__46691),
            .I(N__46566));
    CascadeMux I__10267 (
            .O(N__46690),
            .I(N__46563));
    CascadeMux I__10266 (
            .O(N__46689),
            .I(N__46560));
    CascadeMux I__10265 (
            .O(N__46688),
            .I(N__46557));
    CascadeMux I__10264 (
            .O(N__46687),
            .I(N__46554));
    CascadeMux I__10263 (
            .O(N__46686),
            .I(N__46551));
    CascadeMux I__10262 (
            .O(N__46685),
            .I(N__46548));
    CascadeMux I__10261 (
            .O(N__46684),
            .I(N__46545));
    Span4Mux_v I__10260 (
            .O(N__46681),
            .I(N__46538));
    Span4Mux_h I__10259 (
            .O(N__46678),
            .I(N__46538));
    LocalMux I__10258 (
            .O(N__46669),
            .I(N__46538));
    LocalMux I__10257 (
            .O(N__46664),
            .I(N__46535));
    InMux I__10256 (
            .O(N__46661),
            .I(N__46526));
    InMux I__10255 (
            .O(N__46658),
            .I(N__46526));
    InMux I__10254 (
            .O(N__46655),
            .I(N__46526));
    InMux I__10253 (
            .O(N__46652),
            .I(N__46526));
    InMux I__10252 (
            .O(N__46649),
            .I(N__46517));
    InMux I__10251 (
            .O(N__46646),
            .I(N__46517));
    InMux I__10250 (
            .O(N__46643),
            .I(N__46517));
    InMux I__10249 (
            .O(N__46640),
            .I(N__46517));
    InMux I__10248 (
            .O(N__46637),
            .I(N__46510));
    InMux I__10247 (
            .O(N__46634),
            .I(N__46510));
    InMux I__10246 (
            .O(N__46631),
            .I(N__46510));
    InMux I__10245 (
            .O(N__46628),
            .I(N__46501));
    InMux I__10244 (
            .O(N__46625),
            .I(N__46501));
    InMux I__10243 (
            .O(N__46622),
            .I(N__46501));
    InMux I__10242 (
            .O(N__46619),
            .I(N__46501));
    LocalMux I__10241 (
            .O(N__46610),
            .I(N__46494));
    LocalMux I__10240 (
            .O(N__46601),
            .I(N__46494));
    LocalMux I__10239 (
            .O(N__46592),
            .I(N__46494));
    Span4Mux_v I__10238 (
            .O(N__46587),
            .I(N__46491));
    InMux I__10237 (
            .O(N__46586),
            .I(N__46475));
    InMux I__10236 (
            .O(N__46585),
            .I(N__46468));
    InMux I__10235 (
            .O(N__46584),
            .I(N__46468));
    InMux I__10234 (
            .O(N__46583),
            .I(N__46468));
    InMux I__10233 (
            .O(N__46582),
            .I(N__46459));
    InMux I__10232 (
            .O(N__46581),
            .I(N__46459));
    InMux I__10231 (
            .O(N__46580),
            .I(N__46459));
    InMux I__10230 (
            .O(N__46579),
            .I(N__46459));
    InMux I__10229 (
            .O(N__46578),
            .I(N__46456));
    InMux I__10228 (
            .O(N__46577),
            .I(N__46453));
    InMux I__10227 (
            .O(N__46576),
            .I(N__46450));
    Span12Mux_s11_v I__10226 (
            .O(N__46573),
            .I(N__46439));
    Span4Mux_v I__10225 (
            .O(N__46566),
            .I(N__46436));
    InMux I__10224 (
            .O(N__46563),
            .I(N__46429));
    InMux I__10223 (
            .O(N__46560),
            .I(N__46429));
    InMux I__10222 (
            .O(N__46557),
            .I(N__46429));
    InMux I__10221 (
            .O(N__46554),
            .I(N__46420));
    InMux I__10220 (
            .O(N__46551),
            .I(N__46420));
    InMux I__10219 (
            .O(N__46548),
            .I(N__46420));
    InMux I__10218 (
            .O(N__46545),
            .I(N__46420));
    Span4Mux_v I__10217 (
            .O(N__46538),
            .I(N__46417));
    Span4Mux_v I__10216 (
            .O(N__46535),
            .I(N__46412));
    LocalMux I__10215 (
            .O(N__46526),
            .I(N__46412));
    LocalMux I__10214 (
            .O(N__46517),
            .I(N__46405));
    LocalMux I__10213 (
            .O(N__46510),
            .I(N__46405));
    LocalMux I__10212 (
            .O(N__46501),
            .I(N__46405));
    Span4Mux_v I__10211 (
            .O(N__46494),
            .I(N__46402));
    Sp12to4 I__10210 (
            .O(N__46491),
            .I(N__46399));
    InMux I__10209 (
            .O(N__46490),
            .I(N__46394));
    InMux I__10208 (
            .O(N__46489),
            .I(N__46394));
    CascadeMux I__10207 (
            .O(N__46488),
            .I(N__46390));
    CascadeMux I__10206 (
            .O(N__46487),
            .I(N__46386));
    CascadeMux I__10205 (
            .O(N__46486),
            .I(N__46382));
    CascadeMux I__10204 (
            .O(N__46485),
            .I(N__46377));
    CascadeMux I__10203 (
            .O(N__46484),
            .I(N__46373));
    CascadeMux I__10202 (
            .O(N__46483),
            .I(N__46369));
    CascadeMux I__10201 (
            .O(N__46482),
            .I(N__46365));
    CascadeMux I__10200 (
            .O(N__46481),
            .I(N__46362));
    CascadeMux I__10199 (
            .O(N__46480),
            .I(N__46358));
    CascadeMux I__10198 (
            .O(N__46479),
            .I(N__46354));
    CascadeMux I__10197 (
            .O(N__46478),
            .I(N__46350));
    LocalMux I__10196 (
            .O(N__46475),
            .I(N__46335));
    LocalMux I__10195 (
            .O(N__46468),
            .I(N__46335));
    LocalMux I__10194 (
            .O(N__46459),
            .I(N__46335));
    LocalMux I__10193 (
            .O(N__46456),
            .I(N__46330));
    LocalMux I__10192 (
            .O(N__46453),
            .I(N__46330));
    LocalMux I__10191 (
            .O(N__46450),
            .I(N__46327));
    InMux I__10190 (
            .O(N__46449),
            .I(N__46324));
    InMux I__10189 (
            .O(N__46448),
            .I(N__46317));
    InMux I__10188 (
            .O(N__46447),
            .I(N__46317));
    InMux I__10187 (
            .O(N__46446),
            .I(N__46317));
    InMux I__10186 (
            .O(N__46445),
            .I(N__46308));
    InMux I__10185 (
            .O(N__46444),
            .I(N__46308));
    InMux I__10184 (
            .O(N__46443),
            .I(N__46308));
    InMux I__10183 (
            .O(N__46442),
            .I(N__46308));
    Span12Mux_v I__10182 (
            .O(N__46439),
            .I(N__46301));
    Sp12to4 I__10181 (
            .O(N__46436),
            .I(N__46294));
    LocalMux I__10180 (
            .O(N__46429),
            .I(N__46294));
    LocalMux I__10179 (
            .O(N__46420),
            .I(N__46294));
    Span4Mux_h I__10178 (
            .O(N__46417),
            .I(N__46289));
    Span4Mux_v I__10177 (
            .O(N__46412),
            .I(N__46289));
    Span4Mux_v I__10176 (
            .O(N__46405),
            .I(N__46286));
    Sp12to4 I__10175 (
            .O(N__46402),
            .I(N__46283));
    Span12Mux_h I__10174 (
            .O(N__46399),
            .I(N__46278));
    LocalMux I__10173 (
            .O(N__46394),
            .I(N__46278));
    InMux I__10172 (
            .O(N__46393),
            .I(N__46263));
    InMux I__10171 (
            .O(N__46390),
            .I(N__46263));
    InMux I__10170 (
            .O(N__46389),
            .I(N__46263));
    InMux I__10169 (
            .O(N__46386),
            .I(N__46263));
    InMux I__10168 (
            .O(N__46385),
            .I(N__46263));
    InMux I__10167 (
            .O(N__46382),
            .I(N__46263));
    InMux I__10166 (
            .O(N__46381),
            .I(N__46263));
    InMux I__10165 (
            .O(N__46380),
            .I(N__46246));
    InMux I__10164 (
            .O(N__46377),
            .I(N__46246));
    InMux I__10163 (
            .O(N__46376),
            .I(N__46246));
    InMux I__10162 (
            .O(N__46373),
            .I(N__46246));
    InMux I__10161 (
            .O(N__46372),
            .I(N__46246));
    InMux I__10160 (
            .O(N__46369),
            .I(N__46246));
    InMux I__10159 (
            .O(N__46368),
            .I(N__46246));
    InMux I__10158 (
            .O(N__46365),
            .I(N__46246));
    InMux I__10157 (
            .O(N__46362),
            .I(N__46229));
    InMux I__10156 (
            .O(N__46361),
            .I(N__46229));
    InMux I__10155 (
            .O(N__46358),
            .I(N__46229));
    InMux I__10154 (
            .O(N__46357),
            .I(N__46229));
    InMux I__10153 (
            .O(N__46354),
            .I(N__46229));
    InMux I__10152 (
            .O(N__46353),
            .I(N__46229));
    InMux I__10151 (
            .O(N__46350),
            .I(N__46229));
    InMux I__10150 (
            .O(N__46349),
            .I(N__46229));
    InMux I__10149 (
            .O(N__46348),
            .I(N__46222));
    InMux I__10148 (
            .O(N__46347),
            .I(N__46222));
    InMux I__10147 (
            .O(N__46346),
            .I(N__46222));
    InMux I__10146 (
            .O(N__46345),
            .I(N__46213));
    InMux I__10145 (
            .O(N__46344),
            .I(N__46213));
    InMux I__10144 (
            .O(N__46343),
            .I(N__46213));
    InMux I__10143 (
            .O(N__46342),
            .I(N__46213));
    Span12Mux_v I__10142 (
            .O(N__46335),
            .I(N__46210));
    Span4Mux_v I__10141 (
            .O(N__46330),
            .I(N__46201));
    Span4Mux_v I__10140 (
            .O(N__46327),
            .I(N__46201));
    LocalMux I__10139 (
            .O(N__46324),
            .I(N__46201));
    LocalMux I__10138 (
            .O(N__46317),
            .I(N__46201));
    LocalMux I__10137 (
            .O(N__46308),
            .I(N__46198));
    InMux I__10136 (
            .O(N__46307),
            .I(N__46193));
    InMux I__10135 (
            .O(N__46306),
            .I(N__46193));
    InMux I__10134 (
            .O(N__46305),
            .I(N__46190));
    InMux I__10133 (
            .O(N__46304),
            .I(N__46187));
    Span12Mux_h I__10132 (
            .O(N__46301),
            .I(N__46182));
    Span12Mux_v I__10131 (
            .O(N__46294),
            .I(N__46182));
    Sp12to4 I__10130 (
            .O(N__46289),
            .I(N__46177));
    Sp12to4 I__10129 (
            .O(N__46286),
            .I(N__46177));
    Span12Mux_h I__10128 (
            .O(N__46283),
            .I(N__46162));
    Span12Mux_v I__10127 (
            .O(N__46278),
            .I(N__46162));
    LocalMux I__10126 (
            .O(N__46263),
            .I(N__46162));
    LocalMux I__10125 (
            .O(N__46246),
            .I(N__46162));
    LocalMux I__10124 (
            .O(N__46229),
            .I(N__46162));
    LocalMux I__10123 (
            .O(N__46222),
            .I(N__46162));
    LocalMux I__10122 (
            .O(N__46213),
            .I(N__46162));
    Span12Mux_h I__10121 (
            .O(N__46210),
            .I(N__46159));
    Sp12to4 I__10120 (
            .O(N__46201),
            .I(N__46154));
    Sp12to4 I__10119 (
            .O(N__46198),
            .I(N__46154));
    LocalMux I__10118 (
            .O(N__46193),
            .I(N__46151));
    LocalMux I__10117 (
            .O(N__46190),
            .I(N__46146));
    LocalMux I__10116 (
            .O(N__46187),
            .I(N__46146));
    Span12Mux_h I__10115 (
            .O(N__46182),
            .I(N__46139));
    Span12Mux_h I__10114 (
            .O(N__46177),
            .I(N__46134));
    Span12Mux_v I__10113 (
            .O(N__46162),
            .I(N__46134));
    Span12Mux_h I__10112 (
            .O(N__46159),
            .I(N__46125));
    Span12Mux_v I__10111 (
            .O(N__46154),
            .I(N__46125));
    Sp12to4 I__10110 (
            .O(N__46151),
            .I(N__46125));
    Sp12to4 I__10109 (
            .O(N__46146),
            .I(N__46125));
    InMux I__10108 (
            .O(N__46145),
            .I(N__46122));
    InMux I__10107 (
            .O(N__46144),
            .I(N__46117));
    InMux I__10106 (
            .O(N__46143),
            .I(N__46117));
    InMux I__10105 (
            .O(N__46142),
            .I(N__46114));
    Odrv12 I__10104 (
            .O(N__46139),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10103 (
            .O(N__46134),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10102 (
            .O(N__46125),
            .I(CONSTANT_ONE_NET));
    LocalMux I__10101 (
            .O(N__46122),
            .I(CONSTANT_ONE_NET));
    LocalMux I__10100 (
            .O(N__46117),
            .I(CONSTANT_ONE_NET));
    LocalMux I__10099 (
            .O(N__46114),
            .I(CONSTANT_ONE_NET));
    InMux I__10098 (
            .O(N__46101),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ));
    InMux I__10097 (
            .O(N__46098),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ));
    InMux I__10096 (
            .O(N__46095),
            .I(N__46091));
    InMux I__10095 (
            .O(N__46094),
            .I(N__46088));
    LocalMux I__10094 (
            .O(N__46091),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    LocalMux I__10093 (
            .O(N__46088),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    CascadeMux I__10092 (
            .O(N__46083),
            .I(N__46080));
    InMux I__10091 (
            .O(N__46080),
            .I(N__46077));
    LocalMux I__10090 (
            .O(N__46077),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ));
    InMux I__10089 (
            .O(N__46074),
            .I(N__46070));
    InMux I__10088 (
            .O(N__46073),
            .I(N__46067));
    LocalMux I__10087 (
            .O(N__46070),
            .I(N__46064));
    LocalMux I__10086 (
            .O(N__46067),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__10085 (
            .O(N__46064),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__10084 (
            .O(N__46059),
            .I(N__46056));
    LocalMux I__10083 (
            .O(N__46056),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ));
    InMux I__10082 (
            .O(N__46053),
            .I(N__46049));
    InMux I__10081 (
            .O(N__46052),
            .I(N__46046));
    LocalMux I__10080 (
            .O(N__46049),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_13));
    LocalMux I__10079 (
            .O(N__46046),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_13));
    InMux I__10078 (
            .O(N__46041),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ));
    InMux I__10077 (
            .O(N__46038),
            .I(N__46034));
    InMux I__10076 (
            .O(N__46037),
            .I(N__46031));
    LocalMux I__10075 (
            .O(N__46034),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_14));
    LocalMux I__10074 (
            .O(N__46031),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_14));
    InMux I__10073 (
            .O(N__46026),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ));
    InMux I__10072 (
            .O(N__46023),
            .I(N__46019));
    InMux I__10071 (
            .O(N__46022),
            .I(N__46016));
    LocalMux I__10070 (
            .O(N__46019),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_15));
    LocalMux I__10069 (
            .O(N__46016),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_15));
    InMux I__10068 (
            .O(N__46011),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ));
    InMux I__10067 (
            .O(N__46008),
            .I(bfn_17_10_0_));
    InMux I__10066 (
            .O(N__46005),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ));
    InMux I__10065 (
            .O(N__46002),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ));
    InMux I__10064 (
            .O(N__45999),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ));
    InMux I__10063 (
            .O(N__45996),
            .I(N__45993));
    LocalMux I__10062 (
            .O(N__45993),
            .I(N__45989));
    InMux I__10061 (
            .O(N__45992),
            .I(N__45986));
    Span4Mux_v I__10060 (
            .O(N__45989),
            .I(N__45981));
    LocalMux I__10059 (
            .O(N__45986),
            .I(N__45981));
    Odrv4 I__10058 (
            .O(N__45981),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_20));
    InMux I__10057 (
            .O(N__45978),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ));
    InMux I__10056 (
            .O(N__45975),
            .I(N__45971));
    InMux I__10055 (
            .O(N__45974),
            .I(N__45968));
    LocalMux I__10054 (
            .O(N__45971),
            .I(N__45965));
    LocalMux I__10053 (
            .O(N__45968),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_21));
    Odrv4 I__10052 (
            .O(N__45965),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_21));
    InMux I__10051 (
            .O(N__45960),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ));
    InMux I__10050 (
            .O(N__45957),
            .I(N__45954));
    LocalMux I__10049 (
            .O(N__45954),
            .I(N__45950));
    InMux I__10048 (
            .O(N__45953),
            .I(N__45947));
    Odrv4 I__10047 (
            .O(N__45950),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_5));
    LocalMux I__10046 (
            .O(N__45947),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_5));
    InMux I__10045 (
            .O(N__45942),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ));
    InMux I__10044 (
            .O(N__45939),
            .I(N__45936));
    LocalMux I__10043 (
            .O(N__45936),
            .I(N__45932));
    InMux I__10042 (
            .O(N__45935),
            .I(N__45929));
    Span4Mux_v I__10041 (
            .O(N__45932),
            .I(N__45924));
    LocalMux I__10040 (
            .O(N__45929),
            .I(N__45924));
    Odrv4 I__10039 (
            .O(N__45924),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_6));
    InMux I__10038 (
            .O(N__45921),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ));
    InMux I__10037 (
            .O(N__45918),
            .I(N__45915));
    LocalMux I__10036 (
            .O(N__45915),
            .I(N__45911));
    InMux I__10035 (
            .O(N__45914),
            .I(N__45908));
    Odrv4 I__10034 (
            .O(N__45911),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_7));
    LocalMux I__10033 (
            .O(N__45908),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_7));
    InMux I__10032 (
            .O(N__45903),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ));
    InMux I__10031 (
            .O(N__45900),
            .I(N__45897));
    LocalMux I__10030 (
            .O(N__45897),
            .I(N__45893));
    InMux I__10029 (
            .O(N__45896),
            .I(N__45890));
    Odrv4 I__10028 (
            .O(N__45893),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_8));
    LocalMux I__10027 (
            .O(N__45890),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_8));
    InMux I__10026 (
            .O(N__45885),
            .I(bfn_17_9_0_));
    InMux I__10025 (
            .O(N__45882),
            .I(N__45878));
    InMux I__10024 (
            .O(N__45881),
            .I(N__45875));
    LocalMux I__10023 (
            .O(N__45878),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_9));
    LocalMux I__10022 (
            .O(N__45875),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_9));
    InMux I__10021 (
            .O(N__45870),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ));
    InMux I__10020 (
            .O(N__45867),
            .I(N__45863));
    InMux I__10019 (
            .O(N__45866),
            .I(N__45860));
    LocalMux I__10018 (
            .O(N__45863),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_10));
    LocalMux I__10017 (
            .O(N__45860),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_10));
    InMux I__10016 (
            .O(N__45855),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ));
    InMux I__10015 (
            .O(N__45852),
            .I(N__45848));
    InMux I__10014 (
            .O(N__45851),
            .I(N__45845));
    LocalMux I__10013 (
            .O(N__45848),
            .I(N__45842));
    LocalMux I__10012 (
            .O(N__45845),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_11));
    Odrv4 I__10011 (
            .O(N__45842),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_11));
    InMux I__10010 (
            .O(N__45837),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ));
    InMux I__10009 (
            .O(N__45834),
            .I(N__45831));
    LocalMux I__10008 (
            .O(N__45831),
            .I(N__45827));
    InMux I__10007 (
            .O(N__45830),
            .I(N__45824));
    Odrv4 I__10006 (
            .O(N__45827),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_12));
    LocalMux I__10005 (
            .O(N__45824),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_12));
    InMux I__10004 (
            .O(N__45819),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ));
    InMux I__10003 (
            .O(N__45816),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__10002 (
            .O(N__45813),
            .I(N__45810));
    LocalMux I__10001 (
            .O(N__45810),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__10000 (
            .O(N__45807),
            .I(N__45804));
    LocalMux I__9999 (
            .O(N__45804),
            .I(N__45801));
    Odrv12 I__9998 (
            .O(N__45801),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__9997 (
            .O(N__45798),
            .I(bfn_16_30_0_));
    IoInMux I__9996 (
            .O(N__45795),
            .I(N__45792));
    LocalMux I__9995 (
            .O(N__45792),
            .I(GB_BUFFER_red_c_g_THRU_CO));
    InMux I__9994 (
            .O(N__45789),
            .I(N__45783));
    InMux I__9993 (
            .O(N__45788),
            .I(N__45783));
    LocalMux I__9992 (
            .O(N__45783),
            .I(N__45780));
    Span4Mux_h I__9991 (
            .O(N__45780),
            .I(N__45777));
    Odrv4 I__9990 (
            .O(N__45777),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ));
    InMux I__9989 (
            .O(N__45774),
            .I(N__45771));
    LocalMux I__9988 (
            .O(N__45771),
            .I(\phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ));
    InMux I__9987 (
            .O(N__45768),
            .I(N__45765));
    LocalMux I__9986 (
            .O(N__45765),
            .I(N__45761));
    InMux I__9985 (
            .O(N__45764),
            .I(N__45758));
    Span4Mux_v I__9984 (
            .O(N__45761),
            .I(N__45753));
    LocalMux I__9983 (
            .O(N__45758),
            .I(N__45753));
    Odrv4 I__9982 (
            .O(N__45753),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_1));
    InMux I__9981 (
            .O(N__45750),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ));
    InMux I__9980 (
            .O(N__45747),
            .I(N__45744));
    LocalMux I__9979 (
            .O(N__45744),
            .I(N__45740));
    InMux I__9978 (
            .O(N__45743),
            .I(N__45737));
    Span4Mux_h I__9977 (
            .O(N__45740),
            .I(N__45734));
    LocalMux I__9976 (
            .O(N__45737),
            .I(N__45731));
    Odrv4 I__9975 (
            .O(N__45734),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_2));
    Odrv4 I__9974 (
            .O(N__45731),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_2));
    InMux I__9973 (
            .O(N__45726),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ));
    InMux I__9972 (
            .O(N__45723),
            .I(N__45719));
    InMux I__9971 (
            .O(N__45722),
            .I(N__45716));
    LocalMux I__9970 (
            .O(N__45719),
            .I(N__45713));
    LocalMux I__9969 (
            .O(N__45716),
            .I(N__45710));
    Odrv4 I__9968 (
            .O(N__45713),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_3));
    Odrv4 I__9967 (
            .O(N__45710),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_3));
    InMux I__9966 (
            .O(N__45705),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ));
    InMux I__9965 (
            .O(N__45702),
            .I(N__45698));
    InMux I__9964 (
            .O(N__45701),
            .I(N__45695));
    LocalMux I__9963 (
            .O(N__45698),
            .I(N__45692));
    LocalMux I__9962 (
            .O(N__45695),
            .I(N__45689));
    Odrv4 I__9961 (
            .O(N__45692),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_4));
    Odrv4 I__9960 (
            .O(N__45689),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_4));
    InMux I__9959 (
            .O(N__45684),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ));
    InMux I__9958 (
            .O(N__45681),
            .I(N__45678));
    LocalMux I__9957 (
            .O(N__45678),
            .I(N__45675));
    Span4Mux_s2_v I__9956 (
            .O(N__45675),
            .I(N__45672));
    Span4Mux_v I__9955 (
            .O(N__45672),
            .I(N__45669));
    Sp12to4 I__9954 (
            .O(N__45669),
            .I(N__45666));
    Span12Mux_h I__9953 (
            .O(N__45666),
            .I(N__45663));
    Odrv12 I__9952 (
            .O(N__45663),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__9951 (
            .O(N__45660),
            .I(N__45657));
    InMux I__9950 (
            .O(N__45657),
            .I(N__45654));
    LocalMux I__9949 (
            .O(N__45654),
            .I(N__45651));
    Span4Mux_v I__9948 (
            .O(N__45651),
            .I(N__45648));
    Sp12to4 I__9947 (
            .O(N__45648),
            .I(N__45645));
    Odrv12 I__9946 (
            .O(N__45645),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__9945 (
            .O(N__45642),
            .I(N__45639));
    LocalMux I__9944 (
            .O(N__45639),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__9943 (
            .O(N__45636),
            .I(bfn_16_29_0_));
    InMux I__9942 (
            .O(N__45633),
            .I(N__45630));
    LocalMux I__9941 (
            .O(N__45630),
            .I(N__45627));
    Span4Mux_v I__9940 (
            .O(N__45627),
            .I(N__45624));
    Span4Mux_h I__9939 (
            .O(N__45624),
            .I(N__45621));
    Sp12to4 I__9938 (
            .O(N__45621),
            .I(N__45618));
    Span12Mux_h I__9937 (
            .O(N__45618),
            .I(N__45615));
    Odrv12 I__9936 (
            .O(N__45615),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    CascadeMux I__9935 (
            .O(N__45612),
            .I(N__45609));
    InMux I__9934 (
            .O(N__45609),
            .I(N__45606));
    LocalMux I__9933 (
            .O(N__45606),
            .I(N__45603));
    Span4Mux_s3_v I__9932 (
            .O(N__45603),
            .I(N__45600));
    Span4Mux_h I__9931 (
            .O(N__45600),
            .I(N__45597));
    Span4Mux_h I__9930 (
            .O(N__45597),
            .I(N__45594));
    Odrv4 I__9929 (
            .O(N__45594),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__9928 (
            .O(N__45591),
            .I(N__45588));
    LocalMux I__9927 (
            .O(N__45588),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__9926 (
            .O(N__45585),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__9925 (
            .O(N__45582),
            .I(N__45579));
    LocalMux I__9924 (
            .O(N__45579),
            .I(N__45576));
    Span4Mux_s2_v I__9923 (
            .O(N__45576),
            .I(N__45573));
    Span4Mux_v I__9922 (
            .O(N__45573),
            .I(N__45570));
    Sp12to4 I__9921 (
            .O(N__45570),
            .I(N__45567));
    Span12Mux_h I__9920 (
            .O(N__45567),
            .I(N__45564));
    Odrv12 I__9919 (
            .O(N__45564),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__9918 (
            .O(N__45561),
            .I(N__45558));
    LocalMux I__9917 (
            .O(N__45558),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__9916 (
            .O(N__45555),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__9915 (
            .O(N__45552),
            .I(N__45549));
    InMux I__9914 (
            .O(N__45549),
            .I(N__45546));
    LocalMux I__9913 (
            .O(N__45546),
            .I(N__45543));
    Sp12to4 I__9912 (
            .O(N__45543),
            .I(N__45540));
    Span12Mux_s6_v I__9911 (
            .O(N__45540),
            .I(N__45537));
    Span12Mux_h I__9910 (
            .O(N__45537),
            .I(N__45534));
    Odrv12 I__9909 (
            .O(N__45534),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__9908 (
            .O(N__45531),
            .I(N__45528));
    LocalMux I__9907 (
            .O(N__45528),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__9906 (
            .O(N__45525),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__9905 (
            .O(N__45522),
            .I(N__45519));
    LocalMux I__9904 (
            .O(N__45519),
            .I(N__45516));
    Span12Mux_s6_v I__9903 (
            .O(N__45516),
            .I(N__45513));
    Span12Mux_h I__9902 (
            .O(N__45513),
            .I(N__45510));
    Odrv12 I__9901 (
            .O(N__45510),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__9900 (
            .O(N__45507),
            .I(N__45504));
    LocalMux I__9899 (
            .O(N__45504),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__9898 (
            .O(N__45501),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__9897 (
            .O(N__45498),
            .I(N__45495));
    InMux I__9896 (
            .O(N__45495),
            .I(N__45492));
    LocalMux I__9895 (
            .O(N__45492),
            .I(N__45489));
    Span12Mux_h I__9894 (
            .O(N__45489),
            .I(N__45486));
    Span12Mux_h I__9893 (
            .O(N__45486),
            .I(N__45483));
    Odrv12 I__9892 (
            .O(N__45483),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__9891 (
            .O(N__45480),
            .I(N__45477));
    LocalMux I__9890 (
            .O(N__45477),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__9889 (
            .O(N__45474),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    InMux I__9888 (
            .O(N__45471),
            .I(N__45468));
    LocalMux I__9887 (
            .O(N__45468),
            .I(N__45465));
    Span4Mux_s2_v I__9886 (
            .O(N__45465),
            .I(N__45462));
    Span4Mux_v I__9885 (
            .O(N__45462),
            .I(N__45459));
    Sp12to4 I__9884 (
            .O(N__45459),
            .I(N__45456));
    Span12Mux_h I__9883 (
            .O(N__45456),
            .I(N__45453));
    Odrv12 I__9882 (
            .O(N__45453),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__9881 (
            .O(N__45450),
            .I(N__45447));
    LocalMux I__9880 (
            .O(N__45447),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__9879 (
            .O(N__45444),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__9878 (
            .O(N__45441),
            .I(N__45435));
    CascadeMux I__9877 (
            .O(N__45440),
            .I(N__45431));
    CascadeMux I__9876 (
            .O(N__45439),
            .I(N__45427));
    CascadeMux I__9875 (
            .O(N__45438),
            .I(N__45423));
    LocalMux I__9874 (
            .O(N__45435),
            .I(N__45420));
    InMux I__9873 (
            .O(N__45434),
            .I(N__45407));
    InMux I__9872 (
            .O(N__45431),
            .I(N__45407));
    InMux I__9871 (
            .O(N__45430),
            .I(N__45407));
    InMux I__9870 (
            .O(N__45427),
            .I(N__45407));
    InMux I__9869 (
            .O(N__45426),
            .I(N__45407));
    InMux I__9868 (
            .O(N__45423),
            .I(N__45407));
    Span4Mux_v I__9867 (
            .O(N__45420),
            .I(N__45401));
    LocalMux I__9866 (
            .O(N__45407),
            .I(N__45401));
    InMux I__9865 (
            .O(N__45406),
            .I(N__45398));
    Span4Mux_s2_v I__9864 (
            .O(N__45401),
            .I(N__45395));
    LocalMux I__9863 (
            .O(N__45398),
            .I(N__45392));
    Span4Mux_h I__9862 (
            .O(N__45395),
            .I(N__45389));
    Span12Mux_h I__9861 (
            .O(N__45392),
            .I(N__45386));
    Span4Mux_h I__9860 (
            .O(N__45389),
            .I(N__45383));
    Odrv12 I__9859 (
            .O(N__45386),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    Odrv4 I__9858 (
            .O(N__45383),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__9857 (
            .O(N__45378),
            .I(N__45375));
    InMux I__9856 (
            .O(N__45375),
            .I(N__45372));
    LocalMux I__9855 (
            .O(N__45372),
            .I(N__45369));
    Span4Mux_v I__9854 (
            .O(N__45369),
            .I(N__45366));
    Odrv4 I__9853 (
            .O(N__45366),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__9852 (
            .O(N__45363),
            .I(N__45360));
    LocalMux I__9851 (
            .O(N__45360),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__9850 (
            .O(N__45357),
            .I(N__45354));
    LocalMux I__9849 (
            .O(N__45354),
            .I(N__45351));
    Span4Mux_h I__9848 (
            .O(N__45351),
            .I(N__45348));
    Sp12to4 I__9847 (
            .O(N__45348),
            .I(N__45345));
    Span12Mux_s7_v I__9846 (
            .O(N__45345),
            .I(N__45342));
    Span12Mux_h I__9845 (
            .O(N__45342),
            .I(N__45339));
    Odrv12 I__9844 (
            .O(N__45339),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__9843 (
            .O(N__45336),
            .I(N__45333));
    InMux I__9842 (
            .O(N__45333),
            .I(N__45330));
    LocalMux I__9841 (
            .O(N__45330),
            .I(N__45327));
    Span4Mux_s3_v I__9840 (
            .O(N__45327),
            .I(N__45324));
    Span4Mux_h I__9839 (
            .O(N__45324),
            .I(N__45321));
    Span4Mux_h I__9838 (
            .O(N__45321),
            .I(N__45318));
    Odrv4 I__9837 (
            .O(N__45318),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__9836 (
            .O(N__45315),
            .I(N__45312));
    InMux I__9835 (
            .O(N__45312),
            .I(N__45309));
    LocalMux I__9834 (
            .O(N__45309),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__9833 (
            .O(N__45306),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__9832 (
            .O(N__45303),
            .I(N__45300));
    LocalMux I__9831 (
            .O(N__45300),
            .I(N__45297));
    Span4Mux_s3_v I__9830 (
            .O(N__45297),
            .I(N__45294));
    Span4Mux_v I__9829 (
            .O(N__45294),
            .I(N__45291));
    Sp12to4 I__9828 (
            .O(N__45291),
            .I(N__45288));
    Span12Mux_h I__9827 (
            .O(N__45288),
            .I(N__45285));
    Odrv12 I__9826 (
            .O(N__45285),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__9825 (
            .O(N__45282),
            .I(N__45279));
    InMux I__9824 (
            .O(N__45279),
            .I(N__45276));
    LocalMux I__9823 (
            .O(N__45276),
            .I(N__45273));
    Span4Mux_s3_v I__9822 (
            .O(N__45273),
            .I(N__45270));
    Span4Mux_h I__9821 (
            .O(N__45270),
            .I(N__45267));
    Span4Mux_h I__9820 (
            .O(N__45267),
            .I(N__45264));
    Odrv4 I__9819 (
            .O(N__45264),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__9818 (
            .O(N__45261),
            .I(N__45258));
    LocalMux I__9817 (
            .O(N__45258),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__9816 (
            .O(N__45255),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__9815 (
            .O(N__45252),
            .I(N__45249));
    LocalMux I__9814 (
            .O(N__45249),
            .I(N__45246));
    Span4Mux_h I__9813 (
            .O(N__45246),
            .I(N__45243));
    Span4Mux_h I__9812 (
            .O(N__45243),
            .I(N__45240));
    Span4Mux_h I__9811 (
            .O(N__45240),
            .I(N__45237));
    Odrv4 I__9810 (
            .O(N__45237),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__9809 (
            .O(N__45234),
            .I(N__45231));
    InMux I__9808 (
            .O(N__45231),
            .I(N__45228));
    LocalMux I__9807 (
            .O(N__45228),
            .I(N__45225));
    Sp12to4 I__9806 (
            .O(N__45225),
            .I(N__45222));
    Span12Mux_s7_v I__9805 (
            .O(N__45222),
            .I(N__45219));
    Span12Mux_h I__9804 (
            .O(N__45219),
            .I(N__45216));
    Odrv12 I__9803 (
            .O(N__45216),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    InMux I__9802 (
            .O(N__45213),
            .I(N__45210));
    LocalMux I__9801 (
            .O(N__45210),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__9800 (
            .O(N__45207),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__9799 (
            .O(N__45204),
            .I(N__45201));
    LocalMux I__9798 (
            .O(N__45201),
            .I(N__45198));
    Span12Mux_s7_v I__9797 (
            .O(N__45198),
            .I(N__45195));
    Span12Mux_h I__9796 (
            .O(N__45195),
            .I(N__45192));
    Odrv12 I__9795 (
            .O(N__45192),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__9794 (
            .O(N__45189),
            .I(N__45186));
    InMux I__9793 (
            .O(N__45186),
            .I(N__45183));
    LocalMux I__9792 (
            .O(N__45183),
            .I(N__45180));
    Span12Mux_h I__9791 (
            .O(N__45180),
            .I(N__45177));
    Odrv12 I__9790 (
            .O(N__45177),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__9789 (
            .O(N__45174),
            .I(N__45171));
    LocalMux I__9788 (
            .O(N__45171),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__9787 (
            .O(N__45168),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__9786 (
            .O(N__45165),
            .I(N__45162));
    LocalMux I__9785 (
            .O(N__45162),
            .I(N__45159));
    Span12Mux_h I__9784 (
            .O(N__45159),
            .I(N__45156));
    Span12Mux_h I__9783 (
            .O(N__45156),
            .I(N__45153));
    Odrv12 I__9782 (
            .O(N__45153),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__9781 (
            .O(N__45150),
            .I(N__45147));
    InMux I__9780 (
            .O(N__45147),
            .I(N__45144));
    LocalMux I__9779 (
            .O(N__45144),
            .I(N__45141));
    Span4Mux_v I__9778 (
            .O(N__45141),
            .I(N__45138));
    Sp12to4 I__9777 (
            .O(N__45138),
            .I(N__45135));
    Odrv12 I__9776 (
            .O(N__45135),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__9775 (
            .O(N__45132),
            .I(N__45129));
    LocalMux I__9774 (
            .O(N__45129),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__9773 (
            .O(N__45126),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__9772 (
            .O(N__45123),
            .I(N__45120));
    LocalMux I__9771 (
            .O(N__45120),
            .I(N__45117));
    Span4Mux_v I__9770 (
            .O(N__45117),
            .I(N__45114));
    Span4Mux_h I__9769 (
            .O(N__45114),
            .I(N__45111));
    Sp12to4 I__9768 (
            .O(N__45111),
            .I(N__45108));
    Span12Mux_h I__9767 (
            .O(N__45108),
            .I(N__45105));
    Odrv12 I__9766 (
            .O(N__45105),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__9765 (
            .O(N__45102),
            .I(N__45099));
    InMux I__9764 (
            .O(N__45099),
            .I(N__45096));
    LocalMux I__9763 (
            .O(N__45096),
            .I(N__45093));
    Span12Mux_s5_v I__9762 (
            .O(N__45093),
            .I(N__45090));
    Odrv12 I__9761 (
            .O(N__45090),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__9760 (
            .O(N__45087),
            .I(N__45084));
    LocalMux I__9759 (
            .O(N__45084),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__9758 (
            .O(N__45081),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__9757 (
            .O(N__45078),
            .I(N__45075));
    LocalMux I__9756 (
            .O(N__45075),
            .I(N__45072));
    Span4Mux_h I__9755 (
            .O(N__45072),
            .I(N__45069));
    Span4Mux_h I__9754 (
            .O(N__45069),
            .I(N__45066));
    Sp12to4 I__9753 (
            .O(N__45066),
            .I(N__45063));
    Span12Mux_s7_v I__9752 (
            .O(N__45063),
            .I(N__45060));
    Odrv12 I__9751 (
            .O(N__45060),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__9750 (
            .O(N__45057),
            .I(N__45054));
    InMux I__9749 (
            .O(N__45054),
            .I(N__45051));
    LocalMux I__9748 (
            .O(N__45051),
            .I(N__45048));
    Span4Mux_v I__9747 (
            .O(N__45048),
            .I(N__45045));
    Sp12to4 I__9746 (
            .O(N__45045),
            .I(N__45042));
    Odrv12 I__9745 (
            .O(N__45042),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    InMux I__9744 (
            .O(N__45039),
            .I(N__45036));
    LocalMux I__9743 (
            .O(N__45036),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__9742 (
            .O(N__45033),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    CascadeMux I__9741 (
            .O(N__45030),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ));
    InMux I__9740 (
            .O(N__45027),
            .I(N__45023));
    InMux I__9739 (
            .O(N__45026),
            .I(N__45020));
    LocalMux I__9738 (
            .O(N__45023),
            .I(N__45015));
    LocalMux I__9737 (
            .O(N__45020),
            .I(N__45015));
    Odrv4 I__9736 (
            .O(N__45015),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__9735 (
            .O(N__45012),
            .I(N__45008));
    InMux I__9734 (
            .O(N__45011),
            .I(N__45005));
    LocalMux I__9733 (
            .O(N__45008),
            .I(N__45002));
    LocalMux I__9732 (
            .O(N__45005),
            .I(N__44999));
    Span4Mux_v I__9731 (
            .O(N__45002),
            .I(N__44996));
    Span4Mux_v I__9730 (
            .O(N__44999),
            .I(N__44993));
    Sp12to4 I__9729 (
            .O(N__44996),
            .I(N__44990));
    Span4Mux_h I__9728 (
            .O(N__44993),
            .I(N__44987));
    Span12Mux_h I__9727 (
            .O(N__44990),
            .I(N__44982));
    Sp12to4 I__9726 (
            .O(N__44987),
            .I(N__44982));
    Odrv12 I__9725 (
            .O(N__44982),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    CascadeMux I__9724 (
            .O(N__44979),
            .I(N__44976));
    InMux I__9723 (
            .O(N__44976),
            .I(N__44973));
    LocalMux I__9722 (
            .O(N__44973),
            .I(N__44950));
    InMux I__9721 (
            .O(N__44972),
            .I(N__44944));
    InMux I__9720 (
            .O(N__44971),
            .I(N__44944));
    InMux I__9719 (
            .O(N__44970),
            .I(N__44937));
    InMux I__9718 (
            .O(N__44969),
            .I(N__44937));
    InMux I__9717 (
            .O(N__44968),
            .I(N__44937));
    InMux I__9716 (
            .O(N__44967),
            .I(N__44920));
    InMux I__9715 (
            .O(N__44966),
            .I(N__44920));
    InMux I__9714 (
            .O(N__44965),
            .I(N__44920));
    InMux I__9713 (
            .O(N__44964),
            .I(N__44920));
    InMux I__9712 (
            .O(N__44963),
            .I(N__44920));
    InMux I__9711 (
            .O(N__44962),
            .I(N__44920));
    InMux I__9710 (
            .O(N__44961),
            .I(N__44920));
    InMux I__9709 (
            .O(N__44960),
            .I(N__44920));
    InMux I__9708 (
            .O(N__44959),
            .I(N__44905));
    InMux I__9707 (
            .O(N__44958),
            .I(N__44905));
    InMux I__9706 (
            .O(N__44957),
            .I(N__44905));
    InMux I__9705 (
            .O(N__44956),
            .I(N__44905));
    InMux I__9704 (
            .O(N__44955),
            .I(N__44905));
    InMux I__9703 (
            .O(N__44954),
            .I(N__44905));
    InMux I__9702 (
            .O(N__44953),
            .I(N__44905));
    Span4Mux_v I__9701 (
            .O(N__44950),
            .I(N__44902));
    InMux I__9700 (
            .O(N__44949),
            .I(N__44899));
    LocalMux I__9699 (
            .O(N__44944),
            .I(N__44894));
    LocalMux I__9698 (
            .O(N__44937),
            .I(N__44894));
    LocalMux I__9697 (
            .O(N__44920),
            .I(N__44889));
    LocalMux I__9696 (
            .O(N__44905),
            .I(N__44889));
    Sp12to4 I__9695 (
            .O(N__44902),
            .I(N__44882));
    LocalMux I__9694 (
            .O(N__44899),
            .I(N__44882));
    Span12Mux_s7_v I__9693 (
            .O(N__44894),
            .I(N__44882));
    Span12Mux_s7_h I__9692 (
            .O(N__44889),
            .I(N__44879));
    Span12Mux_h I__9691 (
            .O(N__44882),
            .I(N__44876));
    Odrv12 I__9690 (
            .O(N__44879),
            .I(pwm_duty_input_10));
    Odrv12 I__9689 (
            .O(N__44876),
            .I(pwm_duty_input_10));
    InMux I__9688 (
            .O(N__44871),
            .I(N__44868));
    LocalMux I__9687 (
            .O(N__44868),
            .I(N__44865));
    Span4Mux_v I__9686 (
            .O(N__44865),
            .I(N__44862));
    Sp12to4 I__9685 (
            .O(N__44862),
            .I(N__44859));
    Span12Mux_h I__9684 (
            .O(N__44859),
            .I(N__44856));
    Odrv12 I__9683 (
            .O(N__44856),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__9682 (
            .O(N__44853),
            .I(N__44847));
    InMux I__9681 (
            .O(N__44852),
            .I(N__44847));
    LocalMux I__9680 (
            .O(N__44847),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    CascadeMux I__9679 (
            .O(N__44844),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17_cascade_ ));
    CascadeMux I__9678 (
            .O(N__44841),
            .I(N__44838));
    InMux I__9677 (
            .O(N__44838),
            .I(N__44835));
    LocalMux I__9676 (
            .O(N__44835),
            .I(N__44831));
    InMux I__9675 (
            .O(N__44834),
            .I(N__44828));
    Odrv4 I__9674 (
            .O(N__44831),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    LocalMux I__9673 (
            .O(N__44828),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__9672 (
            .O(N__44823),
            .I(N__44820));
    LocalMux I__9671 (
            .O(N__44820),
            .I(N__44817));
    Span4Mux_s3_v I__9670 (
            .O(N__44817),
            .I(N__44814));
    Span4Mux_v I__9669 (
            .O(N__44814),
            .I(N__44811));
    Sp12to4 I__9668 (
            .O(N__44811),
            .I(N__44808));
    Span12Mux_h I__9667 (
            .O(N__44808),
            .I(N__44805));
    Odrv12 I__9666 (
            .O(N__44805),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__9665 (
            .O(N__44802),
            .I(N__44799));
    InMux I__9664 (
            .O(N__44799),
            .I(N__44796));
    LocalMux I__9663 (
            .O(N__44796),
            .I(N__44793));
    Span4Mux_v I__9662 (
            .O(N__44793),
            .I(N__44790));
    Sp12to4 I__9661 (
            .O(N__44790),
            .I(N__44787));
    Odrv12 I__9660 (
            .O(N__44787),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__9659 (
            .O(N__44784),
            .I(N__44781));
    LocalMux I__9658 (
            .O(N__44781),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__9657 (
            .O(N__44778),
            .I(bfn_16_24_0_));
    InMux I__9656 (
            .O(N__44775),
            .I(\pwm_generator_inst.counter_cry_8 ));
    CascadeMux I__9655 (
            .O(N__44772),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__9654 (
            .O(N__44769),
            .I(N__44766));
    LocalMux I__9653 (
            .O(N__44766),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__9652 (
            .O(N__44763),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__9651 (
            .O(N__44760),
            .I(N__44742));
    InMux I__9650 (
            .O(N__44759),
            .I(N__44742));
    InMux I__9649 (
            .O(N__44758),
            .I(N__44742));
    InMux I__9648 (
            .O(N__44757),
            .I(N__44742));
    InMux I__9647 (
            .O(N__44756),
            .I(N__44733));
    InMux I__9646 (
            .O(N__44755),
            .I(N__44733));
    InMux I__9645 (
            .O(N__44754),
            .I(N__44733));
    InMux I__9644 (
            .O(N__44753),
            .I(N__44733));
    InMux I__9643 (
            .O(N__44752),
            .I(N__44728));
    InMux I__9642 (
            .O(N__44751),
            .I(N__44728));
    LocalMux I__9641 (
            .O(N__44742),
            .I(N__44723));
    LocalMux I__9640 (
            .O(N__44733),
            .I(N__44723));
    LocalMux I__9639 (
            .O(N__44728),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__9638 (
            .O(N__44723),
            .I(\pwm_generator_inst.un1_counter_0 ));
    CascadeMux I__9637 (
            .O(N__44718),
            .I(N__44715));
    InMux I__9636 (
            .O(N__44715),
            .I(N__44712));
    LocalMux I__9635 (
            .O(N__44712),
            .I(N__44708));
    InMux I__9634 (
            .O(N__44711),
            .I(N__44705));
    Odrv4 I__9633 (
            .O(N__44708),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    LocalMux I__9632 (
            .O(N__44705),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__9631 (
            .O(N__44700),
            .I(N__44694));
    InMux I__9630 (
            .O(N__44699),
            .I(N__44694));
    LocalMux I__9629 (
            .O(N__44694),
            .I(N__44691));
    Odrv12 I__9628 (
            .O(N__44691),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__9627 (
            .O(N__44688),
            .I(N__44682));
    InMux I__9626 (
            .O(N__44687),
            .I(N__44682));
    LocalMux I__9625 (
            .O(N__44682),
            .I(N__44679));
    Span4Mux_h I__9624 (
            .O(N__44679),
            .I(N__44676));
    Odrv4 I__9623 (
            .O(N__44676),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    CascadeMux I__9622 (
            .O(N__44673),
            .I(N__44670));
    InMux I__9621 (
            .O(N__44670),
            .I(N__44664));
    InMux I__9620 (
            .O(N__44669),
            .I(N__44664));
    LocalMux I__9619 (
            .O(N__44664),
            .I(N__44661));
    Span4Mux_h I__9618 (
            .O(N__44661),
            .I(N__44658));
    Odrv4 I__9617 (
            .O(N__44658),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__9616 (
            .O(N__44655),
            .I(N__44652));
    LocalMux I__9615 (
            .O(N__44652),
            .I(N__44649));
    Span4Mux_v I__9614 (
            .O(N__44649),
            .I(N__44645));
    InMux I__9613 (
            .O(N__44648),
            .I(N__44642));
    Sp12to4 I__9612 (
            .O(N__44645),
            .I(N__44637));
    LocalMux I__9611 (
            .O(N__44642),
            .I(N__44637));
    Odrv12 I__9610 (
            .O(N__44637),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__9609 (
            .O(N__44634),
            .I(N__44631));
    LocalMux I__9608 (
            .O(N__44631),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__9607 (
            .O(N__44628),
            .I(bfn_16_23_0_));
    InMux I__9606 (
            .O(N__44625),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__9605 (
            .O(N__44622),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__9604 (
            .O(N__44619),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__9603 (
            .O(N__44616),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__9602 (
            .O(N__44613),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__9601 (
            .O(N__44610),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__9600 (
            .O(N__44607),
            .I(\pwm_generator_inst.counter_cry_6 ));
    CascadeMux I__9599 (
            .O(N__44604),
            .I(N__44600));
    InMux I__9598 (
            .O(N__44603),
            .I(N__44597));
    InMux I__9597 (
            .O(N__44600),
            .I(N__44594));
    LocalMux I__9596 (
            .O(N__44597),
            .I(N__44591));
    LocalMux I__9595 (
            .O(N__44594),
            .I(N__44588));
    Span12Mux_s10_v I__9594 (
            .O(N__44591),
            .I(N__44585));
    Span4Mux_h I__9593 (
            .O(N__44588),
            .I(N__44582));
    Odrv12 I__9592 (
            .O(N__44585),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    Odrv4 I__9591 (
            .O(N__44582),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__9590 (
            .O(N__44577),
            .I(N__44571));
    InMux I__9589 (
            .O(N__44576),
            .I(N__44571));
    LocalMux I__9588 (
            .O(N__44571),
            .I(N__44568));
    Odrv12 I__9587 (
            .O(N__44568),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__9586 (
            .O(N__44565),
            .I(N__44559));
    InMux I__9585 (
            .O(N__44564),
            .I(N__44559));
    LocalMux I__9584 (
            .O(N__44559),
            .I(N__44556));
    Odrv12 I__9583 (
            .O(N__44556),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__9582 (
            .O(N__44553),
            .I(N__44549));
    InMux I__9581 (
            .O(N__44552),
            .I(N__44546));
    LocalMux I__9580 (
            .O(N__44549),
            .I(N__44541));
    LocalMux I__9579 (
            .O(N__44546),
            .I(N__44541));
    Odrv12 I__9578 (
            .O(N__44541),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    CascadeMux I__9577 (
            .O(N__44538),
            .I(N__44535));
    InMux I__9576 (
            .O(N__44535),
            .I(N__44532));
    LocalMux I__9575 (
            .O(N__44532),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__9574 (
            .O(N__44529),
            .I(N__44523));
    InMux I__9573 (
            .O(N__44528),
            .I(N__44523));
    LocalMux I__9572 (
            .O(N__44523),
            .I(N__44520));
    Span4Mux_h I__9571 (
            .O(N__44520),
            .I(N__44517));
    Odrv4 I__9570 (
            .O(N__44517),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__9569 (
            .O(N__44514),
            .I(N__44511));
    LocalMux I__9568 (
            .O(N__44511),
            .I(N__44507));
    CascadeMux I__9567 (
            .O(N__44510),
            .I(N__44504));
    Span4Mux_v I__9566 (
            .O(N__44507),
            .I(N__44501));
    InMux I__9565 (
            .O(N__44504),
            .I(N__44498));
    Sp12to4 I__9564 (
            .O(N__44501),
            .I(N__44493));
    LocalMux I__9563 (
            .O(N__44498),
            .I(N__44493));
    Odrv12 I__9562 (
            .O(N__44493),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    CascadeMux I__9561 (
            .O(N__44490),
            .I(N__44487));
    InMux I__9560 (
            .O(N__44487),
            .I(N__44481));
    InMux I__9559 (
            .O(N__44486),
            .I(N__44481));
    LocalMux I__9558 (
            .O(N__44481),
            .I(N__44478));
    Odrv12 I__9557 (
            .O(N__44478),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__9556 (
            .O(N__44475),
            .I(N__44472));
    LocalMux I__9555 (
            .O(N__44472),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    InMux I__9554 (
            .O(N__44469),
            .I(N__44466));
    LocalMux I__9553 (
            .O(N__44466),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__9552 (
            .O(N__44463),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ));
    InMux I__9551 (
            .O(N__44460),
            .I(N__44457));
    LocalMux I__9550 (
            .O(N__44457),
            .I(N__44454));
    Span4Mux_v I__9549 (
            .O(N__44454),
            .I(N__44451));
    Odrv4 I__9548 (
            .O(N__44451),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__9547 (
            .O(N__44448),
            .I(N__44445));
    LocalMux I__9546 (
            .O(N__44445),
            .I(N__44441));
    InMux I__9545 (
            .O(N__44444),
            .I(N__44438));
    Span4Mux_h I__9544 (
            .O(N__44441),
            .I(N__44432));
    LocalMux I__9543 (
            .O(N__44438),
            .I(N__44432));
    InMux I__9542 (
            .O(N__44437),
            .I(N__44429));
    Span4Mux_v I__9541 (
            .O(N__44432),
            .I(N__44425));
    LocalMux I__9540 (
            .O(N__44429),
            .I(N__44422));
    InMux I__9539 (
            .O(N__44428),
            .I(N__44419));
    Sp12to4 I__9538 (
            .O(N__44425),
            .I(N__44414));
    Sp12to4 I__9537 (
            .O(N__44422),
            .I(N__44414));
    LocalMux I__9536 (
            .O(N__44419),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__9535 (
            .O(N__44414),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__9534 (
            .O(N__44409),
            .I(N__44406));
    LocalMux I__9533 (
            .O(N__44406),
            .I(N__44403));
    Span4Mux_v I__9532 (
            .O(N__44403),
            .I(N__44399));
    InMux I__9531 (
            .O(N__44402),
            .I(N__44396));
    Sp12to4 I__9530 (
            .O(N__44399),
            .I(N__44391));
    LocalMux I__9529 (
            .O(N__44396),
            .I(N__44391));
    Odrv12 I__9528 (
            .O(N__44391),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    CascadeMux I__9527 (
            .O(N__44388),
            .I(N__44384));
    InMux I__9526 (
            .O(N__44387),
            .I(N__44381));
    InMux I__9525 (
            .O(N__44384),
            .I(N__44378));
    LocalMux I__9524 (
            .O(N__44381),
            .I(N__44375));
    LocalMux I__9523 (
            .O(N__44378),
            .I(N__44372));
    Span4Mux_h I__9522 (
            .O(N__44375),
            .I(N__44369));
    Span12Mux_h I__9521 (
            .O(N__44372),
            .I(N__44366));
    Span4Mux_h I__9520 (
            .O(N__44369),
            .I(N__44363));
    Odrv12 I__9519 (
            .O(N__44366),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    Odrv4 I__9518 (
            .O(N__44363),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    CascadeMux I__9517 (
            .O(N__44358),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__9516 (
            .O(N__44355),
            .I(N__44352));
    LocalMux I__9515 (
            .O(N__44352),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__9514 (
            .O(N__44349),
            .I(N__44345));
    InMux I__9513 (
            .O(N__44348),
            .I(N__44342));
    LocalMux I__9512 (
            .O(N__44345),
            .I(N__44339));
    LocalMux I__9511 (
            .O(N__44342),
            .I(N__44336));
    Span4Mux_h I__9510 (
            .O(N__44339),
            .I(N__44332));
    Span4Mux_v I__9509 (
            .O(N__44336),
            .I(N__44329));
    InMux I__9508 (
            .O(N__44335),
            .I(N__44326));
    Span4Mux_h I__9507 (
            .O(N__44332),
            .I(N__44323));
    Span4Mux_h I__9506 (
            .O(N__44329),
            .I(N__44320));
    LocalMux I__9505 (
            .O(N__44326),
            .I(N__44317));
    Span4Mux_h I__9504 (
            .O(N__44323),
            .I(N__44314));
    Span4Mux_h I__9503 (
            .O(N__44320),
            .I(N__44311));
    Span4Mux_h I__9502 (
            .O(N__44317),
            .I(N__44306));
    Span4Mux_v I__9501 (
            .O(N__44314),
            .I(N__44306));
    Odrv4 I__9500 (
            .O(N__44311),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__9499 (
            .O(N__44306),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__9498 (
            .O(N__44301),
            .I(N__44298));
    LocalMux I__9497 (
            .O(N__44298),
            .I(N__44295));
    Span4Mux_h I__9496 (
            .O(N__44295),
            .I(N__44292));
    Span4Mux_v I__9495 (
            .O(N__44292),
            .I(N__44288));
    InMux I__9494 (
            .O(N__44291),
            .I(N__44285));
    Odrv4 I__9493 (
            .O(N__44288),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__9492 (
            .O(N__44285),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__9491 (
            .O(N__44280),
            .I(N__44276));
    InMux I__9490 (
            .O(N__44279),
            .I(N__44273));
    LocalMux I__9489 (
            .O(N__44276),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__9488 (
            .O(N__44273),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__9487 (
            .O(N__44268),
            .I(N__44265));
    LocalMux I__9486 (
            .O(N__44265),
            .I(N__44261));
    InMux I__9485 (
            .O(N__44264),
            .I(N__44258));
    Span4Mux_h I__9484 (
            .O(N__44261),
            .I(N__44255));
    LocalMux I__9483 (
            .O(N__44258),
            .I(N__44252));
    Span4Mux_v I__9482 (
            .O(N__44255),
            .I(N__44249));
    Span4Mux_v I__9481 (
            .O(N__44252),
            .I(N__44246));
    Odrv4 I__9480 (
            .O(N__44249),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__9479 (
            .O(N__44246),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__9478 (
            .O(N__44241),
            .I(N__44237));
    InMux I__9477 (
            .O(N__44240),
            .I(N__44234));
    LocalMux I__9476 (
            .O(N__44237),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__9475 (
            .O(N__44234),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__9474 (
            .O(N__44229),
            .I(N__44225));
    InMux I__9473 (
            .O(N__44228),
            .I(N__44222));
    LocalMux I__9472 (
            .O(N__44225),
            .I(N__44219));
    LocalMux I__9471 (
            .O(N__44222),
            .I(N__44216));
    Span4Mux_v I__9470 (
            .O(N__44219),
            .I(N__44213));
    Span4Mux_v I__9469 (
            .O(N__44216),
            .I(N__44208));
    Span4Mux_h I__9468 (
            .O(N__44213),
            .I(N__44208));
    Odrv4 I__9467 (
            .O(N__44208),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    CascadeMux I__9466 (
            .O(N__44205),
            .I(N__44202));
    InMux I__9465 (
            .O(N__44202),
            .I(N__44198));
    InMux I__9464 (
            .O(N__44201),
            .I(N__44195));
    LocalMux I__9463 (
            .O(N__44198),
            .I(N__44192));
    LocalMux I__9462 (
            .O(N__44195),
            .I(N__44189));
    Span4Mux_v I__9461 (
            .O(N__44192),
            .I(N__44184));
    Span4Mux_h I__9460 (
            .O(N__44189),
            .I(N__44184));
    Odrv4 I__9459 (
            .O(N__44184),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    CascadeMux I__9458 (
            .O(N__44181),
            .I(N__44178));
    InMux I__9457 (
            .O(N__44178),
            .I(N__44174));
    InMux I__9456 (
            .O(N__44177),
            .I(N__44171));
    LocalMux I__9455 (
            .O(N__44174),
            .I(N__44168));
    LocalMux I__9454 (
            .O(N__44171),
            .I(N__44165));
    Span4Mux_v I__9453 (
            .O(N__44168),
            .I(N__44162));
    Span4Mux_v I__9452 (
            .O(N__44165),
            .I(N__44157));
    Span4Mux_h I__9451 (
            .O(N__44162),
            .I(N__44157));
    Odrv4 I__9450 (
            .O(N__44157),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__9449 (
            .O(N__44154),
            .I(N__44150));
    InMux I__9448 (
            .O(N__44153),
            .I(N__44147));
    LocalMux I__9447 (
            .O(N__44150),
            .I(N__44144));
    LocalMux I__9446 (
            .O(N__44147),
            .I(N__44141));
    Span4Mux_h I__9445 (
            .O(N__44144),
            .I(N__44138));
    Odrv12 I__9444 (
            .O(N__44141),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    Odrv4 I__9443 (
            .O(N__44138),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__9442 (
            .O(N__44133),
            .I(N__44130));
    LocalMux I__9441 (
            .O(N__44130),
            .I(N__44127));
    Span4Mux_h I__9440 (
            .O(N__44127),
            .I(N__44124));
    Span4Mux_v I__9439 (
            .O(N__44124),
            .I(N__44120));
    InMux I__9438 (
            .O(N__44123),
            .I(N__44117));
    Odrv4 I__9437 (
            .O(N__44120),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    LocalMux I__9436 (
            .O(N__44117),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__9435 (
            .O(N__44112),
            .I(N__44087));
    InMux I__9434 (
            .O(N__44111),
            .I(N__44087));
    InMux I__9433 (
            .O(N__44110),
            .I(N__44078));
    InMux I__9432 (
            .O(N__44109),
            .I(N__44078));
    InMux I__9431 (
            .O(N__44108),
            .I(N__44078));
    InMux I__9430 (
            .O(N__44107),
            .I(N__44078));
    InMux I__9429 (
            .O(N__44106),
            .I(N__44075));
    InMux I__9428 (
            .O(N__44105),
            .I(N__44066));
    InMux I__9427 (
            .O(N__44104),
            .I(N__44061));
    InMux I__9426 (
            .O(N__44103),
            .I(N__44061));
    InMux I__9425 (
            .O(N__44102),
            .I(N__44054));
    InMux I__9424 (
            .O(N__44101),
            .I(N__44054));
    InMux I__9423 (
            .O(N__44100),
            .I(N__44054));
    InMux I__9422 (
            .O(N__44099),
            .I(N__44051));
    InMux I__9421 (
            .O(N__44098),
            .I(N__44048));
    InMux I__9420 (
            .O(N__44097),
            .I(N__44045));
    InMux I__9419 (
            .O(N__44096),
            .I(N__44037));
    InMux I__9418 (
            .O(N__44095),
            .I(N__44037));
    InMux I__9417 (
            .O(N__44094),
            .I(N__44030));
    InMux I__9416 (
            .O(N__44093),
            .I(N__44030));
    InMux I__9415 (
            .O(N__44092),
            .I(N__44030));
    LocalMux I__9414 (
            .O(N__44087),
            .I(N__44023));
    LocalMux I__9413 (
            .O(N__44078),
            .I(N__44023));
    LocalMux I__9412 (
            .O(N__44075),
            .I(N__44023));
    InMux I__9411 (
            .O(N__44074),
            .I(N__44020));
    InMux I__9410 (
            .O(N__44073),
            .I(N__44009));
    InMux I__9409 (
            .O(N__44072),
            .I(N__44009));
    InMux I__9408 (
            .O(N__44071),
            .I(N__44009));
    InMux I__9407 (
            .O(N__44070),
            .I(N__44009));
    InMux I__9406 (
            .O(N__44069),
            .I(N__44009));
    LocalMux I__9405 (
            .O(N__44066),
            .I(N__44002));
    LocalMux I__9404 (
            .O(N__44061),
            .I(N__44002));
    LocalMux I__9403 (
            .O(N__44054),
            .I(N__44002));
    LocalMux I__9402 (
            .O(N__44051),
            .I(N__43995));
    LocalMux I__9401 (
            .O(N__44048),
            .I(N__43995));
    LocalMux I__9400 (
            .O(N__44045),
            .I(N__43995));
    InMux I__9399 (
            .O(N__44044),
            .I(N__43990));
    InMux I__9398 (
            .O(N__44043),
            .I(N__43990));
    InMux I__9397 (
            .O(N__44042),
            .I(N__43987));
    LocalMux I__9396 (
            .O(N__44037),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__9395 (
            .O(N__44030),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__9394 (
            .O(N__44023),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__9393 (
            .O(N__44020),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__9392 (
            .O(N__44009),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__9391 (
            .O(N__44002),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__9390 (
            .O(N__43995),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__9389 (
            .O(N__43990),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__9388 (
            .O(N__43987),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__9387 (
            .O(N__43968),
            .I(N__43964));
    InMux I__9386 (
            .O(N__43967),
            .I(N__43961));
    LocalMux I__9385 (
            .O(N__43964),
            .I(N__43958));
    LocalMux I__9384 (
            .O(N__43961),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    Odrv4 I__9383 (
            .O(N__43958),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    InMux I__9382 (
            .O(N__43953),
            .I(N__43949));
    InMux I__9381 (
            .O(N__43952),
            .I(N__43946));
    LocalMux I__9380 (
            .O(N__43949),
            .I(N__43943));
    LocalMux I__9379 (
            .O(N__43946),
            .I(N__43940));
    Span4Mux_h I__9378 (
            .O(N__43943),
            .I(N__43937));
    Odrv12 I__9377 (
            .O(N__43940),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    Odrv4 I__9376 (
            .O(N__43937),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__9375 (
            .O(N__43932),
            .I(N__43928));
    InMux I__9374 (
            .O(N__43931),
            .I(N__43925));
    LocalMux I__9373 (
            .O(N__43928),
            .I(N__43922));
    LocalMux I__9372 (
            .O(N__43925),
            .I(N__43919));
    Span4Mux_h I__9371 (
            .O(N__43922),
            .I(N__43916));
    Odrv12 I__9370 (
            .O(N__43919),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    Odrv4 I__9369 (
            .O(N__43916),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__9368 (
            .O(N__43911),
            .I(N__43908));
    LocalMux I__9367 (
            .O(N__43908),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__9366 (
            .O(N__43905),
            .I(N__43902));
    LocalMux I__9365 (
            .O(N__43902),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__9364 (
            .O(N__43899),
            .I(N__43896));
    LocalMux I__9363 (
            .O(N__43896),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__9362 (
            .O(N__43893),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ));
    InMux I__9361 (
            .O(N__43890),
            .I(N__43887));
    LocalMux I__9360 (
            .O(N__43887),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    CascadeMux I__9359 (
            .O(N__43884),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ));
    CascadeMux I__9358 (
            .O(N__43881),
            .I(N__43878));
    InMux I__9357 (
            .O(N__43878),
            .I(N__43875));
    LocalMux I__9356 (
            .O(N__43875),
            .I(N__43872));
    Odrv4 I__9355 (
            .O(N__43872),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    InMux I__9354 (
            .O(N__43869),
            .I(N__43866));
    LocalMux I__9353 (
            .O(N__43866),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__9352 (
            .O(N__43863),
            .I(N__43859));
    CascadeMux I__9351 (
            .O(N__43862),
            .I(N__43856));
    LocalMux I__9350 (
            .O(N__43859),
            .I(N__43853));
    InMux I__9349 (
            .O(N__43856),
            .I(N__43850));
    Span4Mux_h I__9348 (
            .O(N__43853),
            .I(N__43845));
    LocalMux I__9347 (
            .O(N__43850),
            .I(N__43845));
    Span4Mux_v I__9346 (
            .O(N__43845),
            .I(N__43842));
    Odrv4 I__9345 (
            .O(N__43842),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__9344 (
            .O(N__43839),
            .I(N__43836));
    LocalMux I__9343 (
            .O(N__43836),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    CascadeMux I__9342 (
            .O(N__43833),
            .I(elapsed_time_ns_1_RNIGF91B_0_4_cascade_));
    InMux I__9341 (
            .O(N__43830),
            .I(N__43827));
    LocalMux I__9340 (
            .O(N__43827),
            .I(N__43824));
    Span4Mux_v I__9339 (
            .O(N__43824),
            .I(N__43821));
    Odrv4 I__9338 (
            .O(N__43821),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ));
    InMux I__9337 (
            .O(N__43818),
            .I(N__43815));
    LocalMux I__9336 (
            .O(N__43815),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    InMux I__9335 (
            .O(N__43812),
            .I(N__43808));
    InMux I__9334 (
            .O(N__43811),
            .I(N__43805));
    LocalMux I__9333 (
            .O(N__43808),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__9332 (
            .O(N__43805),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__9331 (
            .O(N__43800),
            .I(N__43796));
    InMux I__9330 (
            .O(N__43799),
            .I(N__43793));
    LocalMux I__9329 (
            .O(N__43796),
            .I(N__43790));
    LocalMux I__9328 (
            .O(N__43793),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__9327 (
            .O(N__43790),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__9326 (
            .O(N__43785),
            .I(N__43781));
    InMux I__9325 (
            .O(N__43784),
            .I(N__43778));
    LocalMux I__9324 (
            .O(N__43781),
            .I(N__43775));
    LocalMux I__9323 (
            .O(N__43778),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv12 I__9322 (
            .O(N__43775),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__9321 (
            .O(N__43770),
            .I(N__43767));
    LocalMux I__9320 (
            .O(N__43767),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    CascadeMux I__9319 (
            .O(N__43764),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    CascadeMux I__9318 (
            .O(N__43761),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__9317 (
            .O(N__43758),
            .I(N__43755));
    LocalMux I__9316 (
            .O(N__43755),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__9315 (
            .O(N__43752),
            .I(N__43749));
    LocalMux I__9314 (
            .O(N__43749),
            .I(N__43746));
    Span4Mux_h I__9313 (
            .O(N__43746),
            .I(N__43742));
    CascadeMux I__9312 (
            .O(N__43745),
            .I(N__43739));
    Span4Mux_v I__9311 (
            .O(N__43742),
            .I(N__43736));
    InMux I__9310 (
            .O(N__43739),
            .I(N__43733));
    Odrv4 I__9309 (
            .O(N__43736),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__9308 (
            .O(N__43733),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__9307 (
            .O(N__43728),
            .I(N__43725));
    LocalMux I__9306 (
            .O(N__43725),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    CascadeMux I__9305 (
            .O(N__43722),
            .I(elapsed_time_ns_1_RNI2COBB_0_15_cascade_));
    InMux I__9304 (
            .O(N__43719),
            .I(N__43716));
    LocalMux I__9303 (
            .O(N__43716),
            .I(N__43713));
    Span4Mux_v I__9302 (
            .O(N__43713),
            .I(N__43710));
    Odrv4 I__9301 (
            .O(N__43710),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ));
    CascadeMux I__9300 (
            .O(N__43707),
            .I(elapsed_time_ns_1_RNI13CN9_0_14_cascade_));
    InMux I__9299 (
            .O(N__43704),
            .I(N__43698));
    InMux I__9298 (
            .O(N__43703),
            .I(N__43698));
    LocalMux I__9297 (
            .O(N__43698),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__9296 (
            .O(N__43695),
            .I(N__43692));
    LocalMux I__9295 (
            .O(N__43692),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__9294 (
            .O(N__43689),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_));
    InMux I__9293 (
            .O(N__43686),
            .I(N__43683));
    LocalMux I__9292 (
            .O(N__43683),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__9291 (
            .O(N__43680),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    CascadeMux I__9290 (
            .O(N__43677),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__9289 (
            .O(N__43674),
            .I(N__43670));
    InMux I__9288 (
            .O(N__43673),
            .I(N__43667));
    LocalMux I__9287 (
            .O(N__43670),
            .I(N__43664));
    LocalMux I__9286 (
            .O(N__43667),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv12 I__9285 (
            .O(N__43664),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__9284 (
            .O(N__43659),
            .I(N__43655));
    InMux I__9283 (
            .O(N__43658),
            .I(N__43652));
    LocalMux I__9282 (
            .O(N__43655),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__9281 (
            .O(N__43652),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    CascadeMux I__9280 (
            .O(N__43647),
            .I(elapsed_time_ns_1_RNI35CN9_0_16_cascade_));
    InMux I__9279 (
            .O(N__43644),
            .I(N__43641));
    LocalMux I__9278 (
            .O(N__43641),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    CascadeMux I__9277 (
            .O(N__43638),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    InMux I__9276 (
            .O(N__43635),
            .I(N__43632));
    LocalMux I__9275 (
            .O(N__43632),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    CascadeMux I__9274 (
            .O(N__43629),
            .I(elapsed_time_ns_1_RNIG23T9_0_4_cascade_));
    InMux I__9273 (
            .O(N__43626),
            .I(N__43623));
    LocalMux I__9272 (
            .O(N__43623),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    CascadeMux I__9271 (
            .O(N__43620),
            .I(elapsed_time_ns_1_RNI24CN9_0_15_cascade_));
    InMux I__9270 (
            .O(N__43617),
            .I(N__43614));
    LocalMux I__9269 (
            .O(N__43614),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__9268 (
            .O(N__43611),
            .I(N__43608));
    LocalMux I__9267 (
            .O(N__43608),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    CascadeMux I__9266 (
            .O(N__43605),
            .I(elapsed_time_ns_1_RNI57CN9_0_18_cascade_));
    InMux I__9265 (
            .O(N__43602),
            .I(N__43599));
    LocalMux I__9264 (
            .O(N__43599),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    CascadeMux I__9263 (
            .O(N__43596),
            .I(elapsed_time_ns_1_RNIF13T9_0_3_cascade_));
    InMux I__9262 (
            .O(N__43593),
            .I(N__43590));
    LocalMux I__9261 (
            .O(N__43590),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    CascadeMux I__9260 (
            .O(N__43587),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_));
    InMux I__9259 (
            .O(N__43584),
            .I(N__43581));
    LocalMux I__9258 (
            .O(N__43581),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    CascadeMux I__9257 (
            .O(N__43578),
            .I(N__43575));
    InMux I__9256 (
            .O(N__43575),
            .I(N__43569));
    InMux I__9255 (
            .O(N__43574),
            .I(N__43569));
    LocalMux I__9254 (
            .O(N__43569),
            .I(N__43566));
    Span4Mux_v I__9253 (
            .O(N__43566),
            .I(N__43563));
    Odrv4 I__9252 (
            .O(N__43563),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ));
    InMux I__9251 (
            .O(N__43560),
            .I(N__43554));
    InMux I__9250 (
            .O(N__43559),
            .I(N__43554));
    LocalMux I__9249 (
            .O(N__43554),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ));
    InMux I__9248 (
            .O(N__43551),
            .I(N__43548));
    LocalMux I__9247 (
            .O(N__43548),
            .I(N__43545));
    Span4Mux_h I__9246 (
            .O(N__43545),
            .I(N__43542));
    Odrv4 I__9245 (
            .O(N__43542),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ));
    InMux I__9244 (
            .O(N__43539),
            .I(N__43533));
    InMux I__9243 (
            .O(N__43538),
            .I(N__43533));
    LocalMux I__9242 (
            .O(N__43533),
            .I(N__43530));
    Odrv4 I__9241 (
            .O(N__43530),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ));
    InMux I__9240 (
            .O(N__43527),
            .I(N__43521));
    InMux I__9239 (
            .O(N__43526),
            .I(N__43521));
    LocalMux I__9238 (
            .O(N__43521),
            .I(N__43518));
    Odrv4 I__9237 (
            .O(N__43518),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ));
    InMux I__9236 (
            .O(N__43515),
            .I(N__43512));
    LocalMux I__9235 (
            .O(N__43512),
            .I(N__43509));
    Span4Mux_v I__9234 (
            .O(N__43509),
            .I(N__43506));
    Sp12to4 I__9233 (
            .O(N__43506),
            .I(N__43503));
    Odrv12 I__9232 (
            .O(N__43503),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ));
    InMux I__9231 (
            .O(N__43500),
            .I(N__43496));
    InMux I__9230 (
            .O(N__43499),
            .I(N__43493));
    LocalMux I__9229 (
            .O(N__43496),
            .I(N__43490));
    LocalMux I__9228 (
            .O(N__43493),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ));
    Odrv4 I__9227 (
            .O(N__43490),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ));
    InMux I__9226 (
            .O(N__43485),
            .I(N__43481));
    InMux I__9225 (
            .O(N__43484),
            .I(N__43478));
    LocalMux I__9224 (
            .O(N__43481),
            .I(N__43475));
    LocalMux I__9223 (
            .O(N__43478),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ));
    Odrv4 I__9222 (
            .O(N__43475),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ));
    CEMux I__9221 (
            .O(N__43470),
            .I(N__43463));
    CEMux I__9220 (
            .O(N__43469),
            .I(N__43460));
    CEMux I__9219 (
            .O(N__43468),
            .I(N__43457));
    CEMux I__9218 (
            .O(N__43467),
            .I(N__43453));
    CEMux I__9217 (
            .O(N__43466),
            .I(N__43450));
    LocalMux I__9216 (
            .O(N__43463),
            .I(N__43445));
    LocalMux I__9215 (
            .O(N__43460),
            .I(N__43445));
    LocalMux I__9214 (
            .O(N__43457),
            .I(N__43442));
    CEMux I__9213 (
            .O(N__43456),
            .I(N__43439));
    LocalMux I__9212 (
            .O(N__43453),
            .I(N__43436));
    LocalMux I__9211 (
            .O(N__43450),
            .I(N__43432));
    Span4Mux_v I__9210 (
            .O(N__43445),
            .I(N__43425));
    Span4Mux_v I__9209 (
            .O(N__43442),
            .I(N__43425));
    LocalMux I__9208 (
            .O(N__43439),
            .I(N__43425));
    Span4Mux_v I__9207 (
            .O(N__43436),
            .I(N__43422));
    CEMux I__9206 (
            .O(N__43435),
            .I(N__43419));
    Span4Mux_v I__9205 (
            .O(N__43432),
            .I(N__43416));
    Span4Mux_v I__9204 (
            .O(N__43425),
            .I(N__43413));
    Span4Mux_v I__9203 (
            .O(N__43422),
            .I(N__43408));
    LocalMux I__9202 (
            .O(N__43419),
            .I(N__43408));
    Span4Mux_v I__9201 (
            .O(N__43416),
            .I(N__43405));
    Span4Mux_h I__9200 (
            .O(N__43413),
            .I(N__43402));
    Span4Mux_h I__9199 (
            .O(N__43408),
            .I(N__43399));
    Odrv4 I__9198 (
            .O(N__43405),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__9197 (
            .O(N__43402),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__9196 (
            .O(N__43399),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    InMux I__9195 (
            .O(N__43392),
            .I(N__43389));
    LocalMux I__9194 (
            .O(N__43389),
            .I(N__43386));
    Odrv4 I__9193 (
            .O(N__43386),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ));
    InMux I__9192 (
            .O(N__43383),
            .I(N__43380));
    LocalMux I__9191 (
            .O(N__43380),
            .I(N__43377));
    Odrv4 I__9190 (
            .O(N__43377),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ));
    InMux I__9189 (
            .O(N__43374),
            .I(N__43371));
    LocalMux I__9188 (
            .O(N__43371),
            .I(N__43368));
    Span4Mux_h I__9187 (
            .O(N__43368),
            .I(N__43365));
    Odrv4 I__9186 (
            .O(N__43365),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ));
    InMux I__9185 (
            .O(N__43362),
            .I(N__43359));
    LocalMux I__9184 (
            .O(N__43359),
            .I(N__43356));
    Span4Mux_v I__9183 (
            .O(N__43356),
            .I(N__43353));
    Odrv4 I__9182 (
            .O(N__43353),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ));
    InMux I__9181 (
            .O(N__43350),
            .I(N__43347));
    LocalMux I__9180 (
            .O(N__43347),
            .I(N__43344));
    Span4Mux_v I__9179 (
            .O(N__43344),
            .I(N__43341));
    Odrv4 I__9178 (
            .O(N__43341),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ));
    InMux I__9177 (
            .O(N__43338),
            .I(N__43335));
    LocalMux I__9176 (
            .O(N__43335),
            .I(N__43332));
    Span4Mux_h I__9175 (
            .O(N__43332),
            .I(N__43329));
    Odrv4 I__9174 (
            .O(N__43329),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ));
    InMux I__9173 (
            .O(N__43326),
            .I(N__43323));
    LocalMux I__9172 (
            .O(N__43323),
            .I(N__43320));
    Span4Mux_h I__9171 (
            .O(N__43320),
            .I(N__43317));
    Odrv4 I__9170 (
            .O(N__43317),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ));
    CascadeMux I__9169 (
            .O(N__43314),
            .I(N__43310));
    InMux I__9168 (
            .O(N__43313),
            .I(N__43305));
    InMux I__9167 (
            .O(N__43310),
            .I(N__43305));
    LocalMux I__9166 (
            .O(N__43305),
            .I(N__43302));
    Span12Mux_h I__9165 (
            .O(N__43302),
            .I(N__43299));
    Odrv12 I__9164 (
            .O(N__43299),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ));
    InMux I__9163 (
            .O(N__43296),
            .I(N__43293));
    LocalMux I__9162 (
            .O(N__43293),
            .I(N__43290));
    Span4Mux_h I__9161 (
            .O(N__43290),
            .I(N__43287));
    Odrv4 I__9160 (
            .O(N__43287),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ));
    InMux I__9159 (
            .O(N__43284),
            .I(N__43281));
    LocalMux I__9158 (
            .O(N__43281),
            .I(N__43278));
    Span4Mux_h I__9157 (
            .O(N__43278),
            .I(N__43275));
    Odrv4 I__9156 (
            .O(N__43275),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ));
    InMux I__9155 (
            .O(N__43272),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__9154 (
            .O(N__43269),
            .I(N__43266));
    LocalMux I__9153 (
            .O(N__43266),
            .I(N__43263));
    Span4Mux_h I__9152 (
            .O(N__43263),
            .I(N__43260));
    Odrv4 I__9151 (
            .O(N__43260),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ));
    InMux I__9150 (
            .O(N__43257),
            .I(N__43254));
    LocalMux I__9149 (
            .O(N__43254),
            .I(N__43251));
    Span4Mux_h I__9148 (
            .O(N__43251),
            .I(N__43248));
    Odrv4 I__9147 (
            .O(N__43248),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ));
    InMux I__9146 (
            .O(N__43245),
            .I(N__43242));
    LocalMux I__9145 (
            .O(N__43242),
            .I(N__43239));
    Odrv4 I__9144 (
            .O(N__43239),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ));
    InMux I__9143 (
            .O(N__43236),
            .I(N__43233));
    LocalMux I__9142 (
            .O(N__43233),
            .I(N__43230));
    Odrv4 I__9141 (
            .O(N__43230),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ));
    InMux I__9140 (
            .O(N__43227),
            .I(N__43224));
    LocalMux I__9139 (
            .O(N__43224),
            .I(N__43221));
    Odrv4 I__9138 (
            .O(N__43221),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ));
    InMux I__9137 (
            .O(N__43218),
            .I(N__43215));
    LocalMux I__9136 (
            .O(N__43215),
            .I(N__43212));
    Odrv4 I__9135 (
            .O(N__43212),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ));
    InMux I__9134 (
            .O(N__43209),
            .I(N__43206));
    LocalMux I__9133 (
            .O(N__43206),
            .I(N__43203));
    Odrv4 I__9132 (
            .O(N__43203),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ));
    InMux I__9131 (
            .O(N__43200),
            .I(N__43197));
    LocalMux I__9130 (
            .O(N__43197),
            .I(N__43194));
    Odrv4 I__9129 (
            .O(N__43194),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ));
    InMux I__9128 (
            .O(N__43191),
            .I(N__43188));
    LocalMux I__9127 (
            .O(N__43188),
            .I(N__43185));
    Span4Mux_v I__9126 (
            .O(N__43185),
            .I(N__43182));
    Sp12to4 I__9125 (
            .O(N__43182),
            .I(N__43179));
    Odrv12 I__9124 (
            .O(N__43179),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__9123 (
            .O(N__43176),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__9122 (
            .O(N__43173),
            .I(N__43170));
    LocalMux I__9121 (
            .O(N__43170),
            .I(N__43167));
    Span12Mux_s6_v I__9120 (
            .O(N__43167),
            .I(N__43164));
    Odrv12 I__9119 (
            .O(N__43164),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__9118 (
            .O(N__43161),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__9117 (
            .O(N__43158),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__9116 (
            .O(N__43155),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__9115 (
            .O(N__43152),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__9114 (
            .O(N__43149),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__9113 (
            .O(N__43146),
            .I(bfn_15_29_0_));
    CascadeMux I__9112 (
            .O(N__43143),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_));
    InMux I__9111 (
            .O(N__43140),
            .I(N__43137));
    LocalMux I__9110 (
            .O(N__43137),
            .I(N__43134));
    Span4Mux_h I__9109 (
            .O(N__43134),
            .I(N__43131));
    Odrv4 I__9108 (
            .O(N__43131),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ));
    InMux I__9107 (
            .O(N__43128),
            .I(N__43125));
    LocalMux I__9106 (
            .O(N__43125),
            .I(N__43122));
    Span4Mux_v I__9105 (
            .O(N__43122),
            .I(N__43118));
    InMux I__9104 (
            .O(N__43121),
            .I(N__43115));
    Odrv4 I__9103 (
            .O(N__43118),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__9102 (
            .O(N__43115),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9101 (
            .O(N__43110),
            .I(N__43107));
    LocalMux I__9100 (
            .O(N__43107),
            .I(N__43104));
    Span4Mux_v I__9099 (
            .O(N__43104),
            .I(N__43101));
    Span4Mux_v I__9098 (
            .O(N__43101),
            .I(N__43097));
    InMux I__9097 (
            .O(N__43100),
            .I(N__43094));
    Odrv4 I__9096 (
            .O(N__43097),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__9095 (
            .O(N__43094),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    CascadeMux I__9094 (
            .O(N__43089),
            .I(N__43085));
    InMux I__9093 (
            .O(N__43088),
            .I(N__43082));
    InMux I__9092 (
            .O(N__43085),
            .I(N__43079));
    LocalMux I__9091 (
            .O(N__43082),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__9090 (
            .O(N__43079),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__9089 (
            .O(N__43074),
            .I(N__43071));
    LocalMux I__9088 (
            .O(N__43071),
            .I(N__43068));
    Span4Mux_h I__9087 (
            .O(N__43068),
            .I(N__43064));
    InMux I__9086 (
            .O(N__43067),
            .I(N__43061));
    Odrv4 I__9085 (
            .O(N__43064),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__9084 (
            .O(N__43061),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9083 (
            .O(N__43056),
            .I(N__43053));
    LocalMux I__9082 (
            .O(N__43053),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    CascadeMux I__9081 (
            .O(N__43050),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ));
    InMux I__9080 (
            .O(N__43047),
            .I(N__43044));
    LocalMux I__9079 (
            .O(N__43044),
            .I(N__43041));
    Odrv12 I__9078 (
            .O(N__43041),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    InMux I__9077 (
            .O(N__43038),
            .I(N__43035));
    LocalMux I__9076 (
            .O(N__43035),
            .I(N__43032));
    Span4Mux_h I__9075 (
            .O(N__43032),
            .I(N__43028));
    InMux I__9074 (
            .O(N__43031),
            .I(N__43025));
    Odrv4 I__9073 (
            .O(N__43028),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__9072 (
            .O(N__43025),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__9071 (
            .O(N__43020),
            .I(N__43017));
    LocalMux I__9070 (
            .O(N__43017),
            .I(N__43014));
    Span4Mux_h I__9069 (
            .O(N__43014),
            .I(N__43010));
    InMux I__9068 (
            .O(N__43013),
            .I(N__43007));
    Odrv4 I__9067 (
            .O(N__43010),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__9066 (
            .O(N__43007),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__9065 (
            .O(N__43002),
            .I(N__42999));
    LocalMux I__9064 (
            .O(N__42999),
            .I(N__42995));
    CascadeMux I__9063 (
            .O(N__42998),
            .I(N__42992));
    Span4Mux_h I__9062 (
            .O(N__42995),
            .I(N__42989));
    InMux I__9061 (
            .O(N__42992),
            .I(N__42986));
    Odrv4 I__9060 (
            .O(N__42989),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__9059 (
            .O(N__42986),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__9058 (
            .O(N__42981),
            .I(N__42978));
    LocalMux I__9057 (
            .O(N__42978),
            .I(N__42975));
    Span4Mux_h I__9056 (
            .O(N__42975),
            .I(N__42971));
    InMux I__9055 (
            .O(N__42974),
            .I(N__42968));
    Odrv4 I__9054 (
            .O(N__42971),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__9053 (
            .O(N__42968),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__9052 (
            .O(N__42963),
            .I(N__42960));
    LocalMux I__9051 (
            .O(N__42960),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__9050 (
            .O(N__42957),
            .I(N__42954));
    LocalMux I__9049 (
            .O(N__42954),
            .I(N__42951));
    Span12Mux_v I__9048 (
            .O(N__42951),
            .I(N__42947));
    InMux I__9047 (
            .O(N__42950),
            .I(N__42944));
    Odrv12 I__9046 (
            .O(N__42947),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__9045 (
            .O(N__42944),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__9044 (
            .O(N__42939),
            .I(N__42936));
    LocalMux I__9043 (
            .O(N__42936),
            .I(N__42932));
    CascadeMux I__9042 (
            .O(N__42935),
            .I(N__42929));
    Span4Mux_v I__9041 (
            .O(N__42932),
            .I(N__42926));
    InMux I__9040 (
            .O(N__42929),
            .I(N__42923));
    Odrv4 I__9039 (
            .O(N__42926),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__9038 (
            .O(N__42923),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__9037 (
            .O(N__42918),
            .I(N__42915));
    LocalMux I__9036 (
            .O(N__42915),
            .I(N__42912));
    Span4Mux_v I__9035 (
            .O(N__42912),
            .I(N__42909));
    Span4Mux_v I__9034 (
            .O(N__42909),
            .I(N__42905));
    InMux I__9033 (
            .O(N__42908),
            .I(N__42902));
    Odrv4 I__9032 (
            .O(N__42905),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__9031 (
            .O(N__42902),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__9030 (
            .O(N__42897),
            .I(N__42894));
    LocalMux I__9029 (
            .O(N__42894),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__9028 (
            .O(N__42891),
            .I(N__42888));
    LocalMux I__9027 (
            .O(N__42888),
            .I(N__42885));
    Span12Mux_h I__9026 (
            .O(N__42885),
            .I(N__42882));
    Odrv12 I__9025 (
            .O(N__42882),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__9024 (
            .O(N__42879),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__9023 (
            .O(N__42876),
            .I(N__42873));
    LocalMux I__9022 (
            .O(N__42873),
            .I(N__42869));
    InMux I__9021 (
            .O(N__42872),
            .I(N__42866));
    Span4Mux_v I__9020 (
            .O(N__42869),
            .I(N__42863));
    LocalMux I__9019 (
            .O(N__42866),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv4 I__9018 (
            .O(N__42863),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__9017 (
            .O(N__42858),
            .I(N__42855));
    LocalMux I__9016 (
            .O(N__42855),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ));
    InMux I__9015 (
            .O(N__42852),
            .I(N__42849));
    LocalMux I__9014 (
            .O(N__42849),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    CascadeMux I__9013 (
            .O(N__42846),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_));
    InMux I__9012 (
            .O(N__42843),
            .I(N__42840));
    LocalMux I__9011 (
            .O(N__42840),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ));
    InMux I__9010 (
            .O(N__42837),
            .I(N__42834));
    LocalMux I__9009 (
            .O(N__42834),
            .I(N__42831));
    Span4Mux_v I__9008 (
            .O(N__42831),
            .I(N__42827));
    InMux I__9007 (
            .O(N__42830),
            .I(N__42824));
    Odrv4 I__9006 (
            .O(N__42827),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    LocalMux I__9005 (
            .O(N__42824),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__9004 (
            .O(N__42819),
            .I(N__42816));
    LocalMux I__9003 (
            .O(N__42816),
            .I(N__42813));
    Span4Mux_v I__9002 (
            .O(N__42813),
            .I(N__42810));
    Odrv4 I__9001 (
            .O(N__42810),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    InMux I__9000 (
            .O(N__42807),
            .I(N__42804));
    LocalMux I__8999 (
            .O(N__42804),
            .I(N__42801));
    Span4Mux_v I__8998 (
            .O(N__42801),
            .I(N__42798));
    Span4Mux_v I__8997 (
            .O(N__42798),
            .I(N__42794));
    InMux I__8996 (
            .O(N__42797),
            .I(N__42791));
    Odrv4 I__8995 (
            .O(N__42794),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__8994 (
            .O(N__42791),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__8993 (
            .O(N__42786),
            .I(N__42783));
    LocalMux I__8992 (
            .O(N__42783),
            .I(N__42780));
    Span4Mux_h I__8991 (
            .O(N__42780),
            .I(N__42776));
    InMux I__8990 (
            .O(N__42779),
            .I(N__42773));
    Odrv4 I__8989 (
            .O(N__42776),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__8988 (
            .O(N__42773),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__8987 (
            .O(N__42768),
            .I(N__42765));
    LocalMux I__8986 (
            .O(N__42765),
            .I(N__42762));
    Span4Mux_v I__8985 (
            .O(N__42762),
            .I(N__42758));
    CascadeMux I__8984 (
            .O(N__42761),
            .I(N__42755));
    Span4Mux_v I__8983 (
            .O(N__42758),
            .I(N__42752));
    InMux I__8982 (
            .O(N__42755),
            .I(N__42749));
    Odrv4 I__8981 (
            .O(N__42752),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__8980 (
            .O(N__42749),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__8979 (
            .O(N__42744),
            .I(N__42741));
    LocalMux I__8978 (
            .O(N__42741),
            .I(N__42738));
    Span4Mux_v I__8977 (
            .O(N__42738),
            .I(N__42735));
    Span4Mux_v I__8976 (
            .O(N__42735),
            .I(N__42731));
    InMux I__8975 (
            .O(N__42734),
            .I(N__42728));
    Odrv4 I__8974 (
            .O(N__42731),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    LocalMux I__8973 (
            .O(N__42728),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__8972 (
            .O(N__42723),
            .I(N__42720));
    LocalMux I__8971 (
            .O(N__42720),
            .I(N__42717));
    Span4Mux_h I__8970 (
            .O(N__42717),
            .I(N__42713));
    InMux I__8969 (
            .O(N__42716),
            .I(N__42710));
    Odrv4 I__8968 (
            .O(N__42713),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__8967 (
            .O(N__42710),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    CascadeMux I__8966 (
            .O(N__42705),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ));
    InMux I__8965 (
            .O(N__42702),
            .I(N__42699));
    LocalMux I__8964 (
            .O(N__42699),
            .I(N__42696));
    Span4Mux_h I__8963 (
            .O(N__42696),
            .I(N__42693));
    Span4Mux_v I__8962 (
            .O(N__42693),
            .I(N__42689));
    InMux I__8961 (
            .O(N__42692),
            .I(N__42686));
    Odrv4 I__8960 (
            .O(N__42689),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__8959 (
            .O(N__42686),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__8958 (
            .O(N__42681),
            .I(N__42678));
    LocalMux I__8957 (
            .O(N__42678),
            .I(N__42675));
    Odrv12 I__8956 (
            .O(N__42675),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    InMux I__8955 (
            .O(N__42672),
            .I(N__42669));
    LocalMux I__8954 (
            .O(N__42669),
            .I(N__42666));
    Span4Mux_h I__8953 (
            .O(N__42666),
            .I(N__42663));
    Sp12to4 I__8952 (
            .O(N__42663),
            .I(N__42659));
    InMux I__8951 (
            .O(N__42662),
            .I(N__42656));
    Odrv12 I__8950 (
            .O(N__42659),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__8949 (
            .O(N__42656),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__8948 (
            .O(N__42651),
            .I(N__42648));
    LocalMux I__8947 (
            .O(N__42648),
            .I(N__42645));
    Span4Mux_h I__8946 (
            .O(N__42645),
            .I(N__42642));
    Span4Mux_v I__8945 (
            .O(N__42642),
            .I(N__42638));
    InMux I__8944 (
            .O(N__42641),
            .I(N__42635));
    Odrv4 I__8943 (
            .O(N__42638),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__8942 (
            .O(N__42635),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__8941 (
            .O(N__42630),
            .I(N__42627));
    LocalMux I__8940 (
            .O(N__42627),
            .I(N__42624));
    Span4Mux_v I__8939 (
            .O(N__42624),
            .I(N__42620));
    InMux I__8938 (
            .O(N__42623),
            .I(N__42617));
    Odrv4 I__8937 (
            .O(N__42620),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__8936 (
            .O(N__42617),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__8935 (
            .O(N__42612),
            .I(N__42609));
    LocalMux I__8934 (
            .O(N__42609),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__8933 (
            .O(N__42606),
            .I(N__42603));
    LocalMux I__8932 (
            .O(N__42603),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    CascadeMux I__8931 (
            .O(N__42600),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_));
    InMux I__8930 (
            .O(N__42597),
            .I(N__42594));
    LocalMux I__8929 (
            .O(N__42594),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ));
    InMux I__8928 (
            .O(N__42591),
            .I(N__42588));
    LocalMux I__8927 (
            .O(N__42588),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    CascadeMux I__8926 (
            .O(N__42585),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_));
    InMux I__8925 (
            .O(N__42582),
            .I(N__42579));
    LocalMux I__8924 (
            .O(N__42579),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ));
    InMux I__8923 (
            .O(N__42576),
            .I(N__42570));
    InMux I__8922 (
            .O(N__42575),
            .I(N__42570));
    LocalMux I__8921 (
            .O(N__42570),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__8920 (
            .O(N__42567),
            .I(N__42564));
    LocalMux I__8919 (
            .O(N__42564),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    CascadeMux I__8918 (
            .O(N__42561),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_));
    InMux I__8917 (
            .O(N__42558),
            .I(N__42555));
    LocalMux I__8916 (
            .O(N__42555),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ));
    InMux I__8915 (
            .O(N__42552),
            .I(N__42549));
    LocalMux I__8914 (
            .O(N__42549),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ));
    CascadeMux I__8913 (
            .O(N__42546),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_));
    InMux I__8912 (
            .O(N__42543),
            .I(N__42540));
    LocalMux I__8911 (
            .O(N__42540),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ));
    InMux I__8910 (
            .O(N__42537),
            .I(N__42534));
    LocalMux I__8909 (
            .O(N__42534),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    CascadeMux I__8908 (
            .O(N__42531),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    InMux I__8907 (
            .O(N__42528),
            .I(N__42525));
    LocalMux I__8906 (
            .O(N__42525),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ));
    InMux I__8905 (
            .O(N__42522),
            .I(N__42518));
    InMux I__8904 (
            .O(N__42521),
            .I(N__42515));
    LocalMux I__8903 (
            .O(N__42518),
            .I(N__42512));
    LocalMux I__8902 (
            .O(N__42515),
            .I(N__42509));
    Odrv4 I__8901 (
            .O(N__42512),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    Odrv12 I__8900 (
            .O(N__42509),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__8899 (
            .O(N__42504),
            .I(N__42500));
    InMux I__8898 (
            .O(N__42503),
            .I(N__42497));
    LocalMux I__8897 (
            .O(N__42500),
            .I(N__42494));
    LocalMux I__8896 (
            .O(N__42497),
            .I(N__42491));
    Span4Mux_h I__8895 (
            .O(N__42494),
            .I(N__42488));
    Odrv4 I__8894 (
            .O(N__42491),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    Odrv4 I__8893 (
            .O(N__42488),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__8892 (
            .O(N__42483),
            .I(N__42480));
    LocalMux I__8891 (
            .O(N__42480),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    CascadeMux I__8890 (
            .O(N__42477),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_));
    InMux I__8889 (
            .O(N__42474),
            .I(N__42471));
    LocalMux I__8888 (
            .O(N__42471),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ));
    InMux I__8887 (
            .O(N__42468),
            .I(N__42465));
    LocalMux I__8886 (
            .O(N__42465),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ));
    InMux I__8885 (
            .O(N__42462),
            .I(N__42459));
    LocalMux I__8884 (
            .O(N__42459),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    CascadeMux I__8883 (
            .O(N__42456),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_));
    InMux I__8882 (
            .O(N__42453),
            .I(N__42450));
    LocalMux I__8881 (
            .O(N__42450),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ));
    CascadeMux I__8880 (
            .O(N__42447),
            .I(N__42444));
    InMux I__8879 (
            .O(N__42444),
            .I(N__42441));
    LocalMux I__8878 (
            .O(N__42441),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ));
    InMux I__8877 (
            .O(N__42438),
            .I(N__42435));
    LocalMux I__8876 (
            .O(N__42435),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    CascadeMux I__8875 (
            .O(N__42432),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_));
    InMux I__8874 (
            .O(N__42429),
            .I(N__42426));
    LocalMux I__8873 (
            .O(N__42426),
            .I(N__42423));
    Span4Mux_v I__8872 (
            .O(N__42423),
            .I(N__42420));
    Odrv4 I__8871 (
            .O(N__42420),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ));
    InMux I__8870 (
            .O(N__42417),
            .I(N__42414));
    LocalMux I__8869 (
            .O(N__42414),
            .I(N__42410));
    InMux I__8868 (
            .O(N__42413),
            .I(N__42407));
    Span4Mux_h I__8867 (
            .O(N__42410),
            .I(N__42404));
    LocalMux I__8866 (
            .O(N__42407),
            .I(N__42399));
    Span4Mux_h I__8865 (
            .O(N__42404),
            .I(N__42396));
    InMux I__8864 (
            .O(N__42403),
            .I(N__42391));
    InMux I__8863 (
            .O(N__42402),
            .I(N__42391));
    Span4Mux_v I__8862 (
            .O(N__42399),
            .I(N__42388));
    Span4Mux_h I__8861 (
            .O(N__42396),
            .I(N__42385));
    LocalMux I__8860 (
            .O(N__42391),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__8859 (
            .O(N__42388),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__8858 (
            .O(N__42385),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__8857 (
            .O(N__42378),
            .I(N__42374));
    InMux I__8856 (
            .O(N__42377),
            .I(N__42371));
    LocalMux I__8855 (
            .O(N__42374),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__8854 (
            .O(N__42371),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__8853 (
            .O(N__42366),
            .I(N__42363));
    LocalMux I__8852 (
            .O(N__42363),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ));
    InMux I__8851 (
            .O(N__42360),
            .I(N__42357));
    LocalMux I__8850 (
            .O(N__42357),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    CascadeMux I__8849 (
            .O(N__42354),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_));
    InMux I__8848 (
            .O(N__42351),
            .I(N__42348));
    LocalMux I__8847 (
            .O(N__42348),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ));
    InMux I__8846 (
            .O(N__42345),
            .I(N__42342));
    LocalMux I__8845 (
            .O(N__42342),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ));
    InMux I__8844 (
            .O(N__42339),
            .I(N__42336));
    LocalMux I__8843 (
            .O(N__42336),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__8842 (
            .O(N__42333),
            .I(N__42330));
    LocalMux I__8841 (
            .O(N__42330),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    CascadeMux I__8840 (
            .O(N__42327),
            .I(elapsed_time_ns_1_RNIJI91B_0_7_cascade_));
    InMux I__8839 (
            .O(N__42324),
            .I(N__42321));
    LocalMux I__8838 (
            .O(N__42321),
            .I(N__42318));
    Odrv4 I__8837 (
            .O(N__42318),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ));
    InMux I__8836 (
            .O(N__42315),
            .I(N__42309));
    InMux I__8835 (
            .O(N__42314),
            .I(N__42309));
    LocalMux I__8834 (
            .O(N__42309),
            .I(N__42306));
    Span4Mux_v I__8833 (
            .O(N__42306),
            .I(N__42303));
    Span4Mux_v I__8832 (
            .O(N__42303),
            .I(N__42300));
    Odrv4 I__8831 (
            .O(N__42300),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__8830 (
            .O(N__42297),
            .I(N__42291));
    InMux I__8829 (
            .O(N__42296),
            .I(N__42288));
    InMux I__8828 (
            .O(N__42295),
            .I(N__42285));
    InMux I__8827 (
            .O(N__42294),
            .I(N__42282));
    LocalMux I__8826 (
            .O(N__42291),
            .I(N__42277));
    LocalMux I__8825 (
            .O(N__42288),
            .I(N__42274));
    LocalMux I__8824 (
            .O(N__42285),
            .I(N__42271));
    LocalMux I__8823 (
            .O(N__42282),
            .I(N__42268));
    InMux I__8822 (
            .O(N__42281),
            .I(N__42265));
    InMux I__8821 (
            .O(N__42280),
            .I(N__42262));
    Span12Mux_v I__8820 (
            .O(N__42277),
            .I(N__42257));
    Span12Mux_v I__8819 (
            .O(N__42274),
            .I(N__42257));
    Span4Mux_h I__8818 (
            .O(N__42271),
            .I(N__42254));
    Span4Mux_v I__8817 (
            .O(N__42268),
            .I(N__42249));
    LocalMux I__8816 (
            .O(N__42265),
            .I(N__42249));
    LocalMux I__8815 (
            .O(N__42262),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv12 I__8814 (
            .O(N__42257),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__8813 (
            .O(N__42254),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__8812 (
            .O(N__42249),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__8811 (
            .O(N__42240),
            .I(N__42237));
    LocalMux I__8810 (
            .O(N__42237),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    InMux I__8809 (
            .O(N__42234),
            .I(N__42231));
    LocalMux I__8808 (
            .O(N__42231),
            .I(N__42227));
    CascadeMux I__8807 (
            .O(N__42230),
            .I(N__42224));
    Span4Mux_h I__8806 (
            .O(N__42227),
            .I(N__42220));
    InMux I__8805 (
            .O(N__42224),
            .I(N__42217));
    InMux I__8804 (
            .O(N__42223),
            .I(N__42214));
    Odrv4 I__8803 (
            .O(N__42220),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__8802 (
            .O(N__42217),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__8801 (
            .O(N__42214),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__8800 (
            .O(N__42207),
            .I(N__42201));
    InMux I__8799 (
            .O(N__42206),
            .I(N__42201));
    LocalMux I__8798 (
            .O(N__42201),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__8797 (
            .O(N__42198),
            .I(N__42194));
    InMux I__8796 (
            .O(N__42197),
            .I(N__42191));
    LocalMux I__8795 (
            .O(N__42194),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__8794 (
            .O(N__42191),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__8793 (
            .O(N__42186),
            .I(N__42183));
    LocalMux I__8792 (
            .O(N__42183),
            .I(N__42179));
    CascadeMux I__8791 (
            .O(N__42182),
            .I(N__42176));
    Span4Mux_h I__8790 (
            .O(N__42179),
            .I(N__42172));
    InMux I__8789 (
            .O(N__42176),
            .I(N__42169));
    InMux I__8788 (
            .O(N__42175),
            .I(N__42166));
    Odrv4 I__8787 (
            .O(N__42172),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8786 (
            .O(N__42169),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8785 (
            .O(N__42166),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    CEMux I__8784 (
            .O(N__42159),
            .I(N__42154));
    CEMux I__8783 (
            .O(N__42158),
            .I(N__42151));
    CEMux I__8782 (
            .O(N__42157),
            .I(N__42148));
    LocalMux I__8781 (
            .O(N__42154),
            .I(N__42144));
    LocalMux I__8780 (
            .O(N__42151),
            .I(N__42139));
    LocalMux I__8779 (
            .O(N__42148),
            .I(N__42139));
    CEMux I__8778 (
            .O(N__42147),
            .I(N__42136));
    Span4Mux_v I__8777 (
            .O(N__42144),
            .I(N__42128));
    Span4Mux_v I__8776 (
            .O(N__42139),
            .I(N__42128));
    LocalMux I__8775 (
            .O(N__42136),
            .I(N__42128));
    CEMux I__8774 (
            .O(N__42135),
            .I(N__42125));
    Span4Mux_v I__8773 (
            .O(N__42128),
            .I(N__42120));
    LocalMux I__8772 (
            .O(N__42125),
            .I(N__42120));
    Span4Mux_v I__8771 (
            .O(N__42120),
            .I(N__42117));
    Odrv4 I__8770 (
            .O(N__42117),
            .I(\delay_measurement_inst.delay_tr_timer.N_157_i ));
    InMux I__8769 (
            .O(N__42114),
            .I(N__42108));
    InMux I__8768 (
            .O(N__42113),
            .I(N__42108));
    LocalMux I__8767 (
            .O(N__42108),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__8766 (
            .O(N__42105),
            .I(N__42101));
    InMux I__8765 (
            .O(N__42104),
            .I(N__42098));
    LocalMux I__8764 (
            .O(N__42101),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    LocalMux I__8763 (
            .O(N__42098),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__8762 (
            .O(N__42093),
            .I(N__42087));
    InMux I__8761 (
            .O(N__42092),
            .I(N__42087));
    LocalMux I__8760 (
            .O(N__42087),
            .I(N__42084));
    Span4Mux_v I__8759 (
            .O(N__42084),
            .I(N__42081));
    Odrv4 I__8758 (
            .O(N__42081),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__8757 (
            .O(N__42078),
            .I(N__42075));
    LocalMux I__8756 (
            .O(N__42075),
            .I(N__42072));
    Span4Mux_v I__8755 (
            .O(N__42072),
            .I(N__42069));
    Odrv4 I__8754 (
            .O(N__42069),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ));
    InMux I__8753 (
            .O(N__42066),
            .I(N__42063));
    LocalMux I__8752 (
            .O(N__42063),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    CascadeMux I__8751 (
            .O(N__42060),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_));
    InMux I__8750 (
            .O(N__42057),
            .I(N__42054));
    LocalMux I__8749 (
            .O(N__42054),
            .I(N__42051));
    Span4Mux_v I__8748 (
            .O(N__42051),
            .I(N__42048));
    Odrv4 I__8747 (
            .O(N__42048),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ));
    InMux I__8746 (
            .O(N__42045),
            .I(N__42041));
    InMux I__8745 (
            .O(N__42044),
            .I(N__42038));
    LocalMux I__8744 (
            .O(N__42041),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__8743 (
            .O(N__42038),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__8742 (
            .O(N__42033),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    CascadeMux I__8741 (
            .O(N__42030),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__8740 (
            .O(N__42027),
            .I(N__42024));
    LocalMux I__8739 (
            .O(N__42024),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    CascadeMux I__8738 (
            .O(N__42021),
            .I(elapsed_time_ns_1_RNIIH91B_0_6_cascade_));
    CascadeMux I__8737 (
            .O(N__42018),
            .I(N__42015));
    InMux I__8736 (
            .O(N__42015),
            .I(N__42012));
    LocalMux I__8735 (
            .O(N__42012),
            .I(N__42009));
    Odrv4 I__8734 (
            .O(N__42009),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ));
    CascadeMux I__8733 (
            .O(N__42006),
            .I(N__42002));
    InMux I__8732 (
            .O(N__42005),
            .I(N__41997));
    InMux I__8731 (
            .O(N__42002),
            .I(N__41997));
    LocalMux I__8730 (
            .O(N__41997),
            .I(N__41994));
    Span4Mux_v I__8729 (
            .O(N__41994),
            .I(N__41991));
    Odrv4 I__8728 (
            .O(N__41991),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__8727 (
            .O(N__41988),
            .I(N__41985));
    LocalMux I__8726 (
            .O(N__41985),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__8725 (
            .O(N__41982),
            .I(elapsed_time_ns_1_RNI68CN9_0_19_cascade_));
    InMux I__8724 (
            .O(N__41979),
            .I(N__41976));
    LocalMux I__8723 (
            .O(N__41976),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    CascadeMux I__8722 (
            .O(N__41973),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_));
    InMux I__8721 (
            .O(N__41970),
            .I(N__41967));
    LocalMux I__8720 (
            .O(N__41967),
            .I(N__41964));
    Span4Mux_h I__8719 (
            .O(N__41964),
            .I(N__41961));
    Span4Mux_v I__8718 (
            .O(N__41961),
            .I(N__41958));
    Odrv4 I__8717 (
            .O(N__41958),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ));
    InMux I__8716 (
            .O(N__41955),
            .I(N__41952));
    LocalMux I__8715 (
            .O(N__41952),
            .I(N__41949));
    Span4Mux_v I__8714 (
            .O(N__41949),
            .I(N__41946));
    Odrv4 I__8713 (
            .O(N__41946),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ));
    InMux I__8712 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__8711 (
            .O(N__41940),
            .I(N__41937));
    Span12Mux_h I__8710 (
            .O(N__41937),
            .I(N__41934));
    Odrv12 I__8709 (
            .O(N__41934),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ));
    InMux I__8708 (
            .O(N__41931),
            .I(N__41927));
    InMux I__8707 (
            .O(N__41930),
            .I(N__41924));
    LocalMux I__8706 (
            .O(N__41927),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__8705 (
            .O(N__41924),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__8704 (
            .O(N__41919),
            .I(N__41916));
    LocalMux I__8703 (
            .O(N__41916),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    CascadeMux I__8702 (
            .O(N__41913),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    CascadeMux I__8701 (
            .O(N__41910),
            .I(elapsed_time_ns_1_RNIK63T9_0_8_cascade_));
    InMux I__8700 (
            .O(N__41907),
            .I(N__41904));
    LocalMux I__8699 (
            .O(N__41904),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__8698 (
            .O(N__41901),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__8697 (
            .O(N__41898),
            .I(N__41895));
    LocalMux I__8696 (
            .O(N__41895),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    CascadeMux I__8695 (
            .O(N__41892),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_));
    InMux I__8694 (
            .O(N__41889),
            .I(N__41886));
    LocalMux I__8693 (
            .O(N__41886),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    CascadeMux I__8692 (
            .O(N__41883),
            .I(elapsed_time_ns_1_RNIL73T9_0_9_cascade_));
    InMux I__8691 (
            .O(N__41880),
            .I(N__41877));
    LocalMux I__8690 (
            .O(N__41877),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    CascadeMux I__8689 (
            .O(N__41874),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_));
    InMux I__8688 (
            .O(N__41871),
            .I(N__41868));
    LocalMux I__8687 (
            .O(N__41868),
            .I(N__41865));
    Span4Mux_v I__8686 (
            .O(N__41865),
            .I(N__41862));
    Odrv4 I__8685 (
            .O(N__41862),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ));
    CascadeMux I__8684 (
            .O(N__41859),
            .I(N__41856));
    InMux I__8683 (
            .O(N__41856),
            .I(N__41853));
    LocalMux I__8682 (
            .O(N__41853),
            .I(N__41850));
    Odrv4 I__8681 (
            .O(N__41850),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ));
    InMux I__8680 (
            .O(N__41847),
            .I(N__41841));
    InMux I__8679 (
            .O(N__41846),
            .I(N__41841));
    LocalMux I__8678 (
            .O(N__41841),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ));
    InMux I__8677 (
            .O(N__41838),
            .I(N__41835));
    LocalMux I__8676 (
            .O(N__41835),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt16 ));
    InMux I__8675 (
            .O(N__41832),
            .I(N__41826));
    InMux I__8674 (
            .O(N__41831),
            .I(N__41826));
    LocalMux I__8673 (
            .O(N__41826),
            .I(N__41822));
    InMux I__8672 (
            .O(N__41825),
            .I(N__41819));
    Span4Mux_v I__8671 (
            .O(N__41822),
            .I(N__41816));
    LocalMux I__8670 (
            .O(N__41819),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ));
    Odrv4 I__8669 (
            .O(N__41816),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ));
    CascadeMux I__8668 (
            .O(N__41811),
            .I(N__41807));
    CascadeMux I__8667 (
            .O(N__41810),
            .I(N__41804));
    InMux I__8666 (
            .O(N__41807),
            .I(N__41799));
    InMux I__8665 (
            .O(N__41804),
            .I(N__41799));
    LocalMux I__8664 (
            .O(N__41799),
            .I(N__41795));
    InMux I__8663 (
            .O(N__41798),
            .I(N__41792));
    Span4Mux_v I__8662 (
            .O(N__41795),
            .I(N__41789));
    LocalMux I__8661 (
            .O(N__41792),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ));
    Odrv4 I__8660 (
            .O(N__41789),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ));
    CascadeMux I__8659 (
            .O(N__41784),
            .I(N__41781));
    InMux I__8658 (
            .O(N__41781),
            .I(N__41778));
    LocalMux I__8657 (
            .O(N__41778),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ));
    InMux I__8656 (
            .O(N__41775),
            .I(N__41769));
    InMux I__8655 (
            .O(N__41774),
            .I(N__41769));
    LocalMux I__8654 (
            .O(N__41769),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ));
    InMux I__8653 (
            .O(N__41766),
            .I(N__41763));
    LocalMux I__8652 (
            .O(N__41763),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt18 ));
    InMux I__8651 (
            .O(N__41760),
            .I(N__41754));
    InMux I__8650 (
            .O(N__41759),
            .I(N__41754));
    LocalMux I__8649 (
            .O(N__41754),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ));
    InMux I__8648 (
            .O(N__41751),
            .I(N__41745));
    InMux I__8647 (
            .O(N__41750),
            .I(N__41745));
    LocalMux I__8646 (
            .O(N__41745),
            .I(N__41741));
    InMux I__8645 (
            .O(N__41744),
            .I(N__41738));
    Span4Mux_v I__8644 (
            .O(N__41741),
            .I(N__41735));
    LocalMux I__8643 (
            .O(N__41738),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__8642 (
            .O(N__41735),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ));
    CascadeMux I__8641 (
            .O(N__41730),
            .I(N__41726));
    CascadeMux I__8640 (
            .O(N__41729),
            .I(N__41723));
    InMux I__8639 (
            .O(N__41726),
            .I(N__41718));
    InMux I__8638 (
            .O(N__41723),
            .I(N__41718));
    LocalMux I__8637 (
            .O(N__41718),
            .I(N__41714));
    InMux I__8636 (
            .O(N__41717),
            .I(N__41711));
    Span4Mux_v I__8635 (
            .O(N__41714),
            .I(N__41708));
    LocalMux I__8634 (
            .O(N__41711),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ));
    Odrv4 I__8633 (
            .O(N__41708),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ));
    CascadeMux I__8632 (
            .O(N__41703),
            .I(N__41700));
    InMux I__8631 (
            .O(N__41700),
            .I(N__41697));
    LocalMux I__8630 (
            .O(N__41697),
            .I(N__41694));
    Odrv4 I__8629 (
            .O(N__41694),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ));
    InMux I__8628 (
            .O(N__41691),
            .I(N__41688));
    LocalMux I__8627 (
            .O(N__41688),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__8626 (
            .O(N__41685),
            .I(N__41679));
    InMux I__8625 (
            .O(N__41684),
            .I(N__41679));
    LocalMux I__8624 (
            .O(N__41679),
            .I(N__41675));
    InMux I__8623 (
            .O(N__41678),
            .I(N__41672));
    Span4Mux_h I__8622 (
            .O(N__41675),
            .I(N__41669));
    LocalMux I__8621 (
            .O(N__41672),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ));
    Odrv4 I__8620 (
            .O(N__41669),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ));
    InMux I__8619 (
            .O(N__41664),
            .I(N__41658));
    InMux I__8618 (
            .O(N__41663),
            .I(N__41658));
    LocalMux I__8617 (
            .O(N__41658),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ));
    CascadeMux I__8616 (
            .O(N__41655),
            .I(N__41651));
    CascadeMux I__8615 (
            .O(N__41654),
            .I(N__41648));
    InMux I__8614 (
            .O(N__41651),
            .I(N__41643));
    InMux I__8613 (
            .O(N__41648),
            .I(N__41643));
    LocalMux I__8612 (
            .O(N__41643),
            .I(N__41639));
    InMux I__8611 (
            .O(N__41642),
            .I(N__41636));
    Span4Mux_h I__8610 (
            .O(N__41639),
            .I(N__41633));
    LocalMux I__8609 (
            .O(N__41636),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ));
    Odrv4 I__8608 (
            .O(N__41633),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ));
    CascadeMux I__8607 (
            .O(N__41628),
            .I(N__41625));
    InMux I__8606 (
            .O(N__41625),
            .I(N__41622));
    LocalMux I__8605 (
            .O(N__41622),
            .I(N__41619));
    Odrv4 I__8604 (
            .O(N__41619),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ));
    InMux I__8603 (
            .O(N__41616),
            .I(N__41613));
    LocalMux I__8602 (
            .O(N__41613),
            .I(N__41609));
    InMux I__8601 (
            .O(N__41612),
            .I(N__41606));
    Span4Mux_h I__8600 (
            .O(N__41609),
            .I(N__41602));
    LocalMux I__8599 (
            .O(N__41606),
            .I(N__41599));
    InMux I__8598 (
            .O(N__41605),
            .I(N__41596));
    Span4Mux_v I__8597 (
            .O(N__41602),
            .I(N__41593));
    Span12Mux_v I__8596 (
            .O(N__41599),
            .I(N__41590));
    LocalMux I__8595 (
            .O(N__41596),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    Odrv4 I__8594 (
            .O(N__41593),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    Odrv12 I__8593 (
            .O(N__41590),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    CascadeMux I__8592 (
            .O(N__41583),
            .I(N__41579));
    CascadeMux I__8591 (
            .O(N__41582),
            .I(N__41576));
    InMux I__8590 (
            .O(N__41579),
            .I(N__41573));
    InMux I__8589 (
            .O(N__41576),
            .I(N__41570));
    LocalMux I__8588 (
            .O(N__41573),
            .I(N__41565));
    LocalMux I__8587 (
            .O(N__41570),
            .I(N__41565));
    Span4Mux_h I__8586 (
            .O(N__41565),
            .I(N__41561));
    InMux I__8585 (
            .O(N__41564),
            .I(N__41558));
    Span4Mux_v I__8584 (
            .O(N__41561),
            .I(N__41555));
    LocalMux I__8583 (
            .O(N__41558),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ));
    Odrv4 I__8582 (
            .O(N__41555),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ));
    CascadeMux I__8581 (
            .O(N__41550),
            .I(N__41547));
    InMux I__8580 (
            .O(N__41547),
            .I(N__41544));
    LocalMux I__8579 (
            .O(N__41544),
            .I(N__41541));
    Span4Mux_v I__8578 (
            .O(N__41541),
            .I(N__41538));
    Odrv4 I__8577 (
            .O(N__41538),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt24 ));
    InMux I__8576 (
            .O(N__41535),
            .I(N__41532));
    LocalMux I__8575 (
            .O(N__41532),
            .I(N__41529));
    Span4Mux_h I__8574 (
            .O(N__41529),
            .I(N__41526));
    Odrv4 I__8573 (
            .O(N__41526),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt20 ));
    InMux I__8572 (
            .O(N__41523),
            .I(N__41517));
    InMux I__8571 (
            .O(N__41522),
            .I(N__41517));
    LocalMux I__8570 (
            .O(N__41517),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ));
    CascadeMux I__8569 (
            .O(N__41514),
            .I(N__41510));
    CascadeMux I__8568 (
            .O(N__41513),
            .I(N__41507));
    InMux I__8567 (
            .O(N__41510),
            .I(N__41502));
    InMux I__8566 (
            .O(N__41507),
            .I(N__41502));
    LocalMux I__8565 (
            .O(N__41502),
            .I(N__41498));
    InMux I__8564 (
            .O(N__41501),
            .I(N__41495));
    Span4Mux_v I__8563 (
            .O(N__41498),
            .I(N__41492));
    LocalMux I__8562 (
            .O(N__41495),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ));
    Odrv4 I__8561 (
            .O(N__41492),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ));
    InMux I__8560 (
            .O(N__41487),
            .I(N__41481));
    InMux I__8559 (
            .O(N__41486),
            .I(N__41481));
    LocalMux I__8558 (
            .O(N__41481),
            .I(N__41477));
    InMux I__8557 (
            .O(N__41480),
            .I(N__41474));
    Span4Mux_v I__8556 (
            .O(N__41477),
            .I(N__41471));
    LocalMux I__8555 (
            .O(N__41474),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ));
    Odrv4 I__8554 (
            .O(N__41471),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ));
    CascadeMux I__8553 (
            .O(N__41466),
            .I(N__41463));
    InMux I__8552 (
            .O(N__41463),
            .I(N__41460));
    LocalMux I__8551 (
            .O(N__41460),
            .I(N__41457));
    Odrv4 I__8550 (
            .O(N__41457),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ));
    InMux I__8549 (
            .O(N__41454),
            .I(N__41451));
    LocalMux I__8548 (
            .O(N__41451),
            .I(N__41448));
    Span4Mux_h I__8547 (
            .O(N__41448),
            .I(N__41445));
    Odrv4 I__8546 (
            .O(N__41445),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt22 ));
    InMux I__8545 (
            .O(N__41442),
            .I(N__41436));
    InMux I__8544 (
            .O(N__41441),
            .I(N__41436));
    LocalMux I__8543 (
            .O(N__41436),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ));
    InMux I__8542 (
            .O(N__41433),
            .I(N__41427));
    InMux I__8541 (
            .O(N__41432),
            .I(N__41427));
    LocalMux I__8540 (
            .O(N__41427),
            .I(N__41423));
    InMux I__8539 (
            .O(N__41426),
            .I(N__41420));
    Span4Mux_v I__8538 (
            .O(N__41423),
            .I(N__41417));
    LocalMux I__8537 (
            .O(N__41420),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ));
    Odrv4 I__8536 (
            .O(N__41417),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ));
    CascadeMux I__8535 (
            .O(N__41412),
            .I(N__41408));
    CascadeMux I__8534 (
            .O(N__41411),
            .I(N__41405));
    InMux I__8533 (
            .O(N__41408),
            .I(N__41400));
    InMux I__8532 (
            .O(N__41405),
            .I(N__41400));
    LocalMux I__8531 (
            .O(N__41400),
            .I(N__41396));
    InMux I__8530 (
            .O(N__41399),
            .I(N__41393));
    Span12Mux_s11_h I__8529 (
            .O(N__41396),
            .I(N__41390));
    LocalMux I__8528 (
            .O(N__41393),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ));
    Odrv12 I__8527 (
            .O(N__41390),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ));
    InMux I__8526 (
            .O(N__41385),
            .I(N__41382));
    LocalMux I__8525 (
            .O(N__41382),
            .I(N__41379));
    Span4Mux_v I__8524 (
            .O(N__41379),
            .I(N__41376));
    Odrv4 I__8523 (
            .O(N__41376),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ));
    InMux I__8522 (
            .O(N__41373),
            .I(N__41370));
    LocalMux I__8521 (
            .O(N__41370),
            .I(N__41367));
    Odrv4 I__8520 (
            .O(N__41367),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ));
    InMux I__8519 (
            .O(N__41364),
            .I(N__41361));
    LocalMux I__8518 (
            .O(N__41361),
            .I(N__41358));
    Span4Mux_v I__8517 (
            .O(N__41358),
            .I(N__41355));
    Odrv4 I__8516 (
            .O(N__41355),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ));
    InMux I__8515 (
            .O(N__41352),
            .I(N__41349));
    LocalMux I__8514 (
            .O(N__41349),
            .I(N__41346));
    Odrv4 I__8513 (
            .O(N__41346),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ));
    CascadeMux I__8512 (
            .O(N__41343),
            .I(N__41340));
    InMux I__8511 (
            .O(N__41340),
            .I(N__41337));
    LocalMux I__8510 (
            .O(N__41337),
            .I(N__41334));
    Odrv12 I__8509 (
            .O(N__41334),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt20 ));
    InMux I__8508 (
            .O(N__41331),
            .I(N__41325));
    InMux I__8507 (
            .O(N__41330),
            .I(N__41325));
    LocalMux I__8506 (
            .O(N__41325),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ));
    InMux I__8505 (
            .O(N__41322),
            .I(N__41316));
    InMux I__8504 (
            .O(N__41321),
            .I(N__41316));
    LocalMux I__8503 (
            .O(N__41316),
            .I(N__41312));
    InMux I__8502 (
            .O(N__41315),
            .I(N__41309));
    Span4Mux_v I__8501 (
            .O(N__41312),
            .I(N__41306));
    LocalMux I__8500 (
            .O(N__41309),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ));
    Odrv4 I__8499 (
            .O(N__41306),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ));
    CascadeMux I__8498 (
            .O(N__41301),
            .I(N__41297));
    CascadeMux I__8497 (
            .O(N__41300),
            .I(N__41294));
    InMux I__8496 (
            .O(N__41297),
            .I(N__41289));
    InMux I__8495 (
            .O(N__41294),
            .I(N__41289));
    LocalMux I__8494 (
            .O(N__41289),
            .I(N__41285));
    InMux I__8493 (
            .O(N__41288),
            .I(N__41282));
    Span4Mux_v I__8492 (
            .O(N__41285),
            .I(N__41279));
    LocalMux I__8491 (
            .O(N__41282),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ));
    Odrv4 I__8490 (
            .O(N__41279),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ));
    InMux I__8489 (
            .O(N__41274),
            .I(N__41271));
    LocalMux I__8488 (
            .O(N__41271),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ));
    InMux I__8487 (
            .O(N__41268),
            .I(N__41262));
    InMux I__8486 (
            .O(N__41267),
            .I(N__41262));
    LocalMux I__8485 (
            .O(N__41262),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ));
    InMux I__8484 (
            .O(N__41259),
            .I(N__41256));
    LocalMux I__8483 (
            .O(N__41256),
            .I(N__41253));
    Odrv4 I__8482 (
            .O(N__41253),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt22 ));
    IoInMux I__8481 (
            .O(N__41250),
            .I(N__41247));
    LocalMux I__8480 (
            .O(N__41247),
            .I(N__41244));
    Span4Mux_s1_v I__8479 (
            .O(N__41244),
            .I(N__41239));
    InMux I__8478 (
            .O(N__41243),
            .I(N__41234));
    InMux I__8477 (
            .O(N__41242),
            .I(N__41234));
    Odrv4 I__8476 (
            .O(N__41239),
            .I(s1_phy_c));
    LocalMux I__8475 (
            .O(N__41234),
            .I(s1_phy_c));
    InMux I__8474 (
            .O(N__41229),
            .I(N__41224));
    InMux I__8473 (
            .O(N__41228),
            .I(N__41219));
    InMux I__8472 (
            .O(N__41227),
            .I(N__41219));
    LocalMux I__8471 (
            .O(N__41224),
            .I(N__41212));
    LocalMux I__8470 (
            .O(N__41219),
            .I(N__41212));
    CascadeMux I__8469 (
            .O(N__41218),
            .I(N__41208));
    InMux I__8468 (
            .O(N__41217),
            .I(N__41205));
    Span4Mux_s3_v I__8467 (
            .O(N__41212),
            .I(N__41202));
    CascadeMux I__8466 (
            .O(N__41211),
            .I(N__41199));
    InMux I__8465 (
            .O(N__41208),
            .I(N__41196));
    LocalMux I__8464 (
            .O(N__41205),
            .I(N__41193));
    Span4Mux_v I__8463 (
            .O(N__41202),
            .I(N__41190));
    InMux I__8462 (
            .O(N__41199),
            .I(N__41187));
    LocalMux I__8461 (
            .O(N__41196),
            .I(N__41182));
    Span4Mux_h I__8460 (
            .O(N__41193),
            .I(N__41182));
    Span4Mux_v I__8459 (
            .O(N__41190),
            .I(N__41179));
    LocalMux I__8458 (
            .O(N__41187),
            .I(state_3));
    Odrv4 I__8457 (
            .O(N__41182),
            .I(state_3));
    Odrv4 I__8456 (
            .O(N__41179),
            .I(state_3));
    CascadeMux I__8455 (
            .O(N__41172),
            .I(N__41166));
    InMux I__8454 (
            .O(N__41171),
            .I(N__41163));
    InMux I__8453 (
            .O(N__41170),
            .I(N__41156));
    InMux I__8452 (
            .O(N__41169),
            .I(N__41156));
    InMux I__8451 (
            .O(N__41166),
            .I(N__41156));
    LocalMux I__8450 (
            .O(N__41163),
            .I(N__41153));
    LocalMux I__8449 (
            .O(N__41156),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__8448 (
            .O(N__41153),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    CascadeMux I__8447 (
            .O(N__41148),
            .I(N__41145));
    InMux I__8446 (
            .O(N__41145),
            .I(N__41142));
    LocalMux I__8445 (
            .O(N__41142),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ));
    CascadeMux I__8444 (
            .O(N__41139),
            .I(N__41136));
    InMux I__8443 (
            .O(N__41136),
            .I(N__41133));
    LocalMux I__8442 (
            .O(N__41133),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ));
    CascadeMux I__8441 (
            .O(N__41130),
            .I(N__41127));
    InMux I__8440 (
            .O(N__41127),
            .I(N__41124));
    LocalMux I__8439 (
            .O(N__41124),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ));
    CascadeMux I__8438 (
            .O(N__41121),
            .I(N__41118));
    InMux I__8437 (
            .O(N__41118),
            .I(N__41115));
    LocalMux I__8436 (
            .O(N__41115),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ));
    CascadeMux I__8435 (
            .O(N__41112),
            .I(N__41109));
    InMux I__8434 (
            .O(N__41109),
            .I(N__41106));
    LocalMux I__8433 (
            .O(N__41106),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ));
    InMux I__8432 (
            .O(N__41103),
            .I(N__41100));
    LocalMux I__8431 (
            .O(N__41100),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ));
    InMux I__8430 (
            .O(N__41097),
            .I(N__41094));
    LocalMux I__8429 (
            .O(N__41094),
            .I(N__41091));
    Span4Mux_v I__8428 (
            .O(N__41091),
            .I(N__41088));
    Odrv4 I__8427 (
            .O(N__41088),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ));
    InMux I__8426 (
            .O(N__41085),
            .I(N__41082));
    LocalMux I__8425 (
            .O(N__41082),
            .I(N__41079));
    Span4Mux_v I__8424 (
            .O(N__41079),
            .I(N__41076));
    Odrv4 I__8423 (
            .O(N__41076),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ));
    CascadeMux I__8422 (
            .O(N__41073),
            .I(N__41070));
    InMux I__8421 (
            .O(N__41070),
            .I(N__41065));
    InMux I__8420 (
            .O(N__41069),
            .I(N__41062));
    InMux I__8419 (
            .O(N__41068),
            .I(N__41059));
    LocalMux I__8418 (
            .O(N__41065),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__8417 (
            .O(N__41062),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__8416 (
            .O(N__41059),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__8415 (
            .O(N__41052),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__8414 (
            .O(N__41049),
            .I(N__41046));
    InMux I__8413 (
            .O(N__41046),
            .I(N__41041));
    InMux I__8412 (
            .O(N__41045),
            .I(N__41038));
    InMux I__8411 (
            .O(N__41044),
            .I(N__41035));
    LocalMux I__8410 (
            .O(N__41041),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__8409 (
            .O(N__41038),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__8408 (
            .O(N__41035),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__8407 (
            .O(N__41028),
            .I(bfn_14_27_0_));
    InMux I__8406 (
            .O(N__41025),
            .I(N__41020));
    InMux I__8405 (
            .O(N__41024),
            .I(N__41017));
    InMux I__8404 (
            .O(N__41023),
            .I(N__41014));
    LocalMux I__8403 (
            .O(N__41020),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__8402 (
            .O(N__41017),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__8401 (
            .O(N__41014),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__8400 (
            .O(N__41007),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8399 (
            .O(N__41004),
            .I(N__41000));
    InMux I__8398 (
            .O(N__41003),
            .I(N__40997));
    LocalMux I__8397 (
            .O(N__41000),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__8396 (
            .O(N__40997),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__8395 (
            .O(N__40992),
            .I(N__40989));
    InMux I__8394 (
            .O(N__40989),
            .I(N__40984));
    InMux I__8393 (
            .O(N__40988),
            .I(N__40981));
    InMux I__8392 (
            .O(N__40987),
            .I(N__40978));
    LocalMux I__8391 (
            .O(N__40984),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__8390 (
            .O(N__40981),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__8389 (
            .O(N__40978),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__8388 (
            .O(N__40971),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__8387 (
            .O(N__40968),
            .I(N__40964));
    InMux I__8386 (
            .O(N__40967),
            .I(N__40961));
    LocalMux I__8385 (
            .O(N__40964),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__8384 (
            .O(N__40961),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__8383 (
            .O(N__40956),
            .I(N__40951));
    CascadeMux I__8382 (
            .O(N__40955),
            .I(N__40948));
    InMux I__8381 (
            .O(N__40954),
            .I(N__40945));
    InMux I__8380 (
            .O(N__40951),
            .I(N__40940));
    InMux I__8379 (
            .O(N__40948),
            .I(N__40940));
    LocalMux I__8378 (
            .O(N__40945),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__8377 (
            .O(N__40940),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__8376 (
            .O(N__40935),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8375 (
            .O(N__40932),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8374 (
            .O(N__40929),
            .I(N__40926));
    LocalMux I__8373 (
            .O(N__40926),
            .I(N__40922));
    InMux I__8372 (
            .O(N__40925),
            .I(N__40918));
    Span4Mux_v I__8371 (
            .O(N__40922),
            .I(N__40915));
    InMux I__8370 (
            .O(N__40921),
            .I(N__40911));
    LocalMux I__8369 (
            .O(N__40918),
            .I(N__40908));
    Span4Mux_h I__8368 (
            .O(N__40915),
            .I(N__40905));
    InMux I__8367 (
            .O(N__40914),
            .I(N__40902));
    LocalMux I__8366 (
            .O(N__40911),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__8365 (
            .O(N__40908),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__8364 (
            .O(N__40905),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__8363 (
            .O(N__40902),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__8362 (
            .O(N__40893),
            .I(N__40888));
    InMux I__8361 (
            .O(N__40892),
            .I(N__40882));
    InMux I__8360 (
            .O(N__40891),
            .I(N__40882));
    LocalMux I__8359 (
            .O(N__40888),
            .I(N__40879));
    InMux I__8358 (
            .O(N__40887),
            .I(N__40876));
    LocalMux I__8357 (
            .O(N__40882),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__8356 (
            .O(N__40879),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__8355 (
            .O(N__40876),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    CascadeMux I__8354 (
            .O(N__40869),
            .I(N__40866));
    InMux I__8353 (
            .O(N__40866),
            .I(N__40861));
    InMux I__8352 (
            .O(N__40865),
            .I(N__40858));
    InMux I__8351 (
            .O(N__40864),
            .I(N__40855));
    LocalMux I__8350 (
            .O(N__40861),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__8349 (
            .O(N__40858),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__8348 (
            .O(N__40855),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__8347 (
            .O(N__40848),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__8346 (
            .O(N__40845),
            .I(N__40842));
    InMux I__8345 (
            .O(N__40842),
            .I(N__40837));
    InMux I__8344 (
            .O(N__40841),
            .I(N__40834));
    InMux I__8343 (
            .O(N__40840),
            .I(N__40831));
    LocalMux I__8342 (
            .O(N__40837),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8341 (
            .O(N__40834),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8340 (
            .O(N__40831),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__8339 (
            .O(N__40824),
            .I(bfn_14_26_0_));
    CascadeMux I__8338 (
            .O(N__40821),
            .I(N__40818));
    InMux I__8337 (
            .O(N__40818),
            .I(N__40813));
    InMux I__8336 (
            .O(N__40817),
            .I(N__40810));
    InMux I__8335 (
            .O(N__40816),
            .I(N__40807));
    LocalMux I__8334 (
            .O(N__40813),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__8333 (
            .O(N__40810),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__8332 (
            .O(N__40807),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__8331 (
            .O(N__40800),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__8330 (
            .O(N__40797),
            .I(N__40792));
    InMux I__8329 (
            .O(N__40796),
            .I(N__40787));
    InMux I__8328 (
            .O(N__40795),
            .I(N__40787));
    LocalMux I__8327 (
            .O(N__40792),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__8326 (
            .O(N__40787),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__8325 (
            .O(N__40782),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__8324 (
            .O(N__40779),
            .I(N__40776));
    InMux I__8323 (
            .O(N__40776),
            .I(N__40771));
    InMux I__8322 (
            .O(N__40775),
            .I(N__40768));
    InMux I__8321 (
            .O(N__40774),
            .I(N__40765));
    LocalMux I__8320 (
            .O(N__40771),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__8319 (
            .O(N__40768),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__8318 (
            .O(N__40765),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__8317 (
            .O(N__40758),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__8316 (
            .O(N__40755),
            .I(N__40750));
    CascadeMux I__8315 (
            .O(N__40754),
            .I(N__40747));
    InMux I__8314 (
            .O(N__40753),
            .I(N__40744));
    InMux I__8313 (
            .O(N__40750),
            .I(N__40739));
    InMux I__8312 (
            .O(N__40747),
            .I(N__40739));
    LocalMux I__8311 (
            .O(N__40744),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__8310 (
            .O(N__40739),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__8309 (
            .O(N__40734),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__8308 (
            .O(N__40731),
            .I(N__40728));
    InMux I__8307 (
            .O(N__40728),
            .I(N__40723));
    InMux I__8306 (
            .O(N__40727),
            .I(N__40720));
    InMux I__8305 (
            .O(N__40726),
            .I(N__40717));
    LocalMux I__8304 (
            .O(N__40723),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__8303 (
            .O(N__40720),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__8302 (
            .O(N__40717),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__8301 (
            .O(N__40710),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__8300 (
            .O(N__40707),
            .I(N__40704));
    InMux I__8299 (
            .O(N__40704),
            .I(N__40699));
    InMux I__8298 (
            .O(N__40703),
            .I(N__40696));
    InMux I__8297 (
            .O(N__40702),
            .I(N__40693));
    LocalMux I__8296 (
            .O(N__40699),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__8295 (
            .O(N__40696),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__8294 (
            .O(N__40693),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__8293 (
            .O(N__40686),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8292 (
            .O(N__40683),
            .I(N__40680));
    InMux I__8291 (
            .O(N__40680),
            .I(N__40675));
    InMux I__8290 (
            .O(N__40679),
            .I(N__40672));
    InMux I__8289 (
            .O(N__40678),
            .I(N__40669));
    LocalMux I__8288 (
            .O(N__40675),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__8287 (
            .O(N__40672),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__8286 (
            .O(N__40669),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__8285 (
            .O(N__40662),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__8284 (
            .O(N__40659),
            .I(N__40656));
    InMux I__8283 (
            .O(N__40656),
            .I(N__40651));
    InMux I__8282 (
            .O(N__40655),
            .I(N__40648));
    InMux I__8281 (
            .O(N__40654),
            .I(N__40645));
    LocalMux I__8280 (
            .O(N__40651),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__8279 (
            .O(N__40648),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__8278 (
            .O(N__40645),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__8277 (
            .O(N__40638),
            .I(bfn_14_25_0_));
    InMux I__8276 (
            .O(N__40635),
            .I(N__40630));
    InMux I__8275 (
            .O(N__40634),
            .I(N__40627));
    InMux I__8274 (
            .O(N__40633),
            .I(N__40624));
    LocalMux I__8273 (
            .O(N__40630),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__8272 (
            .O(N__40627),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__8271 (
            .O(N__40624),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__8270 (
            .O(N__40617),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__8269 (
            .O(N__40614),
            .I(N__40611));
    InMux I__8268 (
            .O(N__40611),
            .I(N__40606));
    InMux I__8267 (
            .O(N__40610),
            .I(N__40603));
    InMux I__8266 (
            .O(N__40609),
            .I(N__40600));
    LocalMux I__8265 (
            .O(N__40606),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__8264 (
            .O(N__40603),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__8263 (
            .O(N__40600),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__8262 (
            .O(N__40593),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__8261 (
            .O(N__40590),
            .I(N__40585));
    CascadeMux I__8260 (
            .O(N__40589),
            .I(N__40582));
    InMux I__8259 (
            .O(N__40588),
            .I(N__40579));
    InMux I__8258 (
            .O(N__40585),
            .I(N__40574));
    InMux I__8257 (
            .O(N__40582),
            .I(N__40574));
    LocalMux I__8256 (
            .O(N__40579),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__8255 (
            .O(N__40574),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__8254 (
            .O(N__40569),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__8253 (
            .O(N__40566),
            .I(N__40563));
    InMux I__8252 (
            .O(N__40563),
            .I(N__40558));
    InMux I__8251 (
            .O(N__40562),
            .I(N__40555));
    InMux I__8250 (
            .O(N__40561),
            .I(N__40552));
    LocalMux I__8249 (
            .O(N__40558),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__8248 (
            .O(N__40555),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__8247 (
            .O(N__40552),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__8246 (
            .O(N__40545),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__8245 (
            .O(N__40542),
            .I(N__40539));
    InMux I__8244 (
            .O(N__40539),
            .I(N__40534));
    InMux I__8243 (
            .O(N__40538),
            .I(N__40531));
    InMux I__8242 (
            .O(N__40537),
            .I(N__40528));
    LocalMux I__8241 (
            .O(N__40534),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__8240 (
            .O(N__40531),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__8239 (
            .O(N__40528),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__8238 (
            .O(N__40521),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__8237 (
            .O(N__40518),
            .I(N__40515));
    InMux I__8236 (
            .O(N__40515),
            .I(N__40510));
    InMux I__8235 (
            .O(N__40514),
            .I(N__40507));
    InMux I__8234 (
            .O(N__40513),
            .I(N__40504));
    LocalMux I__8233 (
            .O(N__40510),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__8232 (
            .O(N__40507),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__8231 (
            .O(N__40504),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__8230 (
            .O(N__40497),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__8229 (
            .O(N__40494),
            .I(N__40490));
    InMux I__8228 (
            .O(N__40493),
            .I(N__40487));
    LocalMux I__8227 (
            .O(N__40490),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ));
    LocalMux I__8226 (
            .O(N__40487),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ));
    InMux I__8225 (
            .O(N__40482),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ));
    InMux I__8224 (
            .O(N__40479),
            .I(N__40476));
    LocalMux I__8223 (
            .O(N__40476),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ));
    InMux I__8222 (
            .O(N__40473),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ));
    InMux I__8221 (
            .O(N__40470),
            .I(N__40467));
    LocalMux I__8220 (
            .O(N__40467),
            .I(N__40464));
    Span12Mux_h I__8219 (
            .O(N__40464),
            .I(N__40460));
    InMux I__8218 (
            .O(N__40463),
            .I(N__40457));
    Span12Mux_v I__8217 (
            .O(N__40460),
            .I(N__40454));
    LocalMux I__8216 (
            .O(N__40457),
            .I(N__40451));
    Odrv12 I__8215 (
            .O(N__40454),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_28));
    Odrv4 I__8214 (
            .O(N__40451),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_28));
    InMux I__8213 (
            .O(N__40446),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__8212 (
            .O(N__40443),
            .I(N__40438));
    InMux I__8211 (
            .O(N__40442),
            .I(N__40433));
    InMux I__8210 (
            .O(N__40441),
            .I(N__40433));
    LocalMux I__8209 (
            .O(N__40438),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__8208 (
            .O(N__40433),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__8207 (
            .O(N__40428),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__8206 (
            .O(N__40425),
            .I(N__40422));
    InMux I__8205 (
            .O(N__40422),
            .I(N__40417));
    InMux I__8204 (
            .O(N__40421),
            .I(N__40414));
    InMux I__8203 (
            .O(N__40420),
            .I(N__40411));
    LocalMux I__8202 (
            .O(N__40417),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__8201 (
            .O(N__40414),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__8200 (
            .O(N__40411),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__8199 (
            .O(N__40404),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__8198 (
            .O(N__40401),
            .I(N__40396));
    CascadeMux I__8197 (
            .O(N__40400),
            .I(N__40393));
    InMux I__8196 (
            .O(N__40399),
            .I(N__40390));
    InMux I__8195 (
            .O(N__40396),
            .I(N__40385));
    InMux I__8194 (
            .O(N__40393),
            .I(N__40385));
    LocalMux I__8193 (
            .O(N__40390),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__8192 (
            .O(N__40385),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__8191 (
            .O(N__40380),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__8190 (
            .O(N__40377),
            .I(N__40374));
    InMux I__8189 (
            .O(N__40374),
            .I(N__40369));
    InMux I__8188 (
            .O(N__40373),
            .I(N__40366));
    InMux I__8187 (
            .O(N__40372),
            .I(N__40363));
    LocalMux I__8186 (
            .O(N__40369),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__8185 (
            .O(N__40366),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__8184 (
            .O(N__40363),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__8183 (
            .O(N__40356),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__8182 (
            .O(N__40353),
            .I(N__40350));
    InMux I__8181 (
            .O(N__40350),
            .I(N__40345));
    InMux I__8180 (
            .O(N__40349),
            .I(N__40342));
    InMux I__8179 (
            .O(N__40348),
            .I(N__40339));
    LocalMux I__8178 (
            .O(N__40345),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__8177 (
            .O(N__40342),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__8176 (
            .O(N__40339),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__8175 (
            .O(N__40332),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__8174 (
            .O(N__40329),
            .I(N__40325));
    InMux I__8173 (
            .O(N__40328),
            .I(N__40322));
    LocalMux I__8172 (
            .O(N__40325),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ));
    LocalMux I__8171 (
            .O(N__40322),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ));
    InMux I__8170 (
            .O(N__40317),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ));
    InMux I__8169 (
            .O(N__40314),
            .I(N__40310));
    InMux I__8168 (
            .O(N__40313),
            .I(N__40307));
    LocalMux I__8167 (
            .O(N__40310),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ));
    LocalMux I__8166 (
            .O(N__40307),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ));
    InMux I__8165 (
            .O(N__40302),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ));
    InMux I__8164 (
            .O(N__40299),
            .I(N__40295));
    InMux I__8163 (
            .O(N__40298),
            .I(N__40292));
    LocalMux I__8162 (
            .O(N__40295),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ));
    LocalMux I__8161 (
            .O(N__40292),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ));
    InMux I__8160 (
            .O(N__40287),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ));
    InMux I__8159 (
            .O(N__40284),
            .I(N__40280));
    InMux I__8158 (
            .O(N__40283),
            .I(N__40277));
    LocalMux I__8157 (
            .O(N__40280),
            .I(N__40274));
    LocalMux I__8156 (
            .O(N__40277),
            .I(N__40271));
    Odrv4 I__8155 (
            .O(N__40274),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ));
    Odrv4 I__8154 (
            .O(N__40271),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ));
    InMux I__8153 (
            .O(N__40266),
            .I(bfn_14_23_0_));
    InMux I__8152 (
            .O(N__40263),
            .I(N__40259));
    InMux I__8151 (
            .O(N__40262),
            .I(N__40256));
    LocalMux I__8150 (
            .O(N__40259),
            .I(N__40251));
    LocalMux I__8149 (
            .O(N__40256),
            .I(N__40251));
    Odrv4 I__8148 (
            .O(N__40251),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ));
    InMux I__8147 (
            .O(N__40248),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ));
    InMux I__8146 (
            .O(N__40245),
            .I(N__40241));
    InMux I__8145 (
            .O(N__40244),
            .I(N__40238));
    LocalMux I__8144 (
            .O(N__40241),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ));
    LocalMux I__8143 (
            .O(N__40238),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ));
    InMux I__8142 (
            .O(N__40233),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ));
    InMux I__8141 (
            .O(N__40230),
            .I(N__40226));
    InMux I__8140 (
            .O(N__40229),
            .I(N__40223));
    LocalMux I__8139 (
            .O(N__40226),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ));
    LocalMux I__8138 (
            .O(N__40223),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ));
    InMux I__8137 (
            .O(N__40218),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ));
    InMux I__8136 (
            .O(N__40215),
            .I(N__40211));
    InMux I__8135 (
            .O(N__40214),
            .I(N__40208));
    LocalMux I__8134 (
            .O(N__40211),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ));
    LocalMux I__8133 (
            .O(N__40208),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ));
    InMux I__8132 (
            .O(N__40203),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ));
    InMux I__8131 (
            .O(N__40200),
            .I(N__40196));
    InMux I__8130 (
            .O(N__40199),
            .I(N__40193));
    LocalMux I__8129 (
            .O(N__40196),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ));
    LocalMux I__8128 (
            .O(N__40193),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ));
    InMux I__8127 (
            .O(N__40188),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ));
    InMux I__8126 (
            .O(N__40185),
            .I(N__40181));
    InMux I__8125 (
            .O(N__40184),
            .I(N__40178));
    LocalMux I__8124 (
            .O(N__40181),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ));
    LocalMux I__8123 (
            .O(N__40178),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ));
    InMux I__8122 (
            .O(N__40173),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ));
    InMux I__8121 (
            .O(N__40170),
            .I(N__40166));
    InMux I__8120 (
            .O(N__40169),
            .I(N__40163));
    LocalMux I__8119 (
            .O(N__40166),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ));
    LocalMux I__8118 (
            .O(N__40163),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ));
    InMux I__8117 (
            .O(N__40158),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ));
    InMux I__8116 (
            .O(N__40155),
            .I(N__40151));
    InMux I__8115 (
            .O(N__40154),
            .I(N__40148));
    LocalMux I__8114 (
            .O(N__40151),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ));
    LocalMux I__8113 (
            .O(N__40148),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ));
    InMux I__8112 (
            .O(N__40143),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ));
    InMux I__8111 (
            .O(N__40140),
            .I(N__40136));
    InMux I__8110 (
            .O(N__40139),
            .I(N__40133));
    LocalMux I__8109 (
            .O(N__40136),
            .I(N__40130));
    LocalMux I__8108 (
            .O(N__40133),
            .I(N__40127));
    Odrv4 I__8107 (
            .O(N__40130),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ));
    Odrv4 I__8106 (
            .O(N__40127),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ));
    InMux I__8105 (
            .O(N__40122),
            .I(bfn_14_22_0_));
    InMux I__8104 (
            .O(N__40119),
            .I(N__40115));
    InMux I__8103 (
            .O(N__40118),
            .I(N__40112));
    LocalMux I__8102 (
            .O(N__40115),
            .I(N__40107));
    LocalMux I__8101 (
            .O(N__40112),
            .I(N__40107));
    Odrv4 I__8100 (
            .O(N__40107),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ));
    InMux I__8099 (
            .O(N__40104),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ));
    InMux I__8098 (
            .O(N__40101),
            .I(N__40097));
    InMux I__8097 (
            .O(N__40100),
            .I(N__40094));
    LocalMux I__8096 (
            .O(N__40097),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ));
    LocalMux I__8095 (
            .O(N__40094),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ));
    InMux I__8094 (
            .O(N__40089),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ));
    InMux I__8093 (
            .O(N__40086),
            .I(N__40083));
    LocalMux I__8092 (
            .O(N__40083),
            .I(N__40079));
    InMux I__8091 (
            .O(N__40082),
            .I(N__40076));
    Span4Mux_h I__8090 (
            .O(N__40079),
            .I(N__40073));
    LocalMux I__8089 (
            .O(N__40076),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ));
    Odrv4 I__8088 (
            .O(N__40073),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ));
    InMux I__8087 (
            .O(N__40068),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ));
    InMux I__8086 (
            .O(N__40065),
            .I(N__40061));
    InMux I__8085 (
            .O(N__40064),
            .I(N__40058));
    LocalMux I__8084 (
            .O(N__40061),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ));
    LocalMux I__8083 (
            .O(N__40058),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ));
    InMux I__8082 (
            .O(N__40053),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ));
    InMux I__8081 (
            .O(N__40050),
            .I(N__40046));
    InMux I__8080 (
            .O(N__40049),
            .I(N__40043));
    LocalMux I__8079 (
            .O(N__40046),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ));
    LocalMux I__8078 (
            .O(N__40043),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ));
    InMux I__8077 (
            .O(N__40038),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ));
    InMux I__8076 (
            .O(N__40035),
            .I(N__40031));
    InMux I__8075 (
            .O(N__40034),
            .I(N__40028));
    LocalMux I__8074 (
            .O(N__40031),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ));
    LocalMux I__8073 (
            .O(N__40028),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ));
    InMux I__8072 (
            .O(N__40023),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ));
    InMux I__8071 (
            .O(N__40020),
            .I(N__40016));
    InMux I__8070 (
            .O(N__40019),
            .I(N__40013));
    LocalMux I__8069 (
            .O(N__40016),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ));
    LocalMux I__8068 (
            .O(N__40013),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ));
    InMux I__8067 (
            .O(N__40008),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ));
    InMux I__8066 (
            .O(N__40005),
            .I(N__40001));
    InMux I__8065 (
            .O(N__40004),
            .I(N__39998));
    LocalMux I__8064 (
            .O(N__40001),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ));
    LocalMux I__8063 (
            .O(N__39998),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ));
    InMux I__8062 (
            .O(N__39993),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ));
    InMux I__8061 (
            .O(N__39990),
            .I(N__39987));
    LocalMux I__8060 (
            .O(N__39987),
            .I(N__39984));
    Span4Mux_v I__8059 (
            .O(N__39984),
            .I(N__39981));
    Odrv4 I__8058 (
            .O(N__39981),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ));
    InMux I__8057 (
            .O(N__39978),
            .I(N__39974));
    InMux I__8056 (
            .O(N__39977),
            .I(N__39971));
    LocalMux I__8055 (
            .O(N__39974),
            .I(N__39968));
    LocalMux I__8054 (
            .O(N__39971),
            .I(N__39965));
    Odrv4 I__8053 (
            .O(N__39968),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ));
    Odrv4 I__8052 (
            .O(N__39965),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ));
    InMux I__8051 (
            .O(N__39960),
            .I(bfn_14_21_0_));
    InMux I__8050 (
            .O(N__39957),
            .I(N__39953));
    InMux I__8049 (
            .O(N__39956),
            .I(N__39950));
    LocalMux I__8048 (
            .O(N__39953),
            .I(N__39945));
    LocalMux I__8047 (
            .O(N__39950),
            .I(N__39945));
    Odrv4 I__8046 (
            .O(N__39945),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ));
    InMux I__8045 (
            .O(N__39942),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ));
    InMux I__8044 (
            .O(N__39939),
            .I(N__39935));
    InMux I__8043 (
            .O(N__39938),
            .I(N__39932));
    LocalMux I__8042 (
            .O(N__39935),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ));
    LocalMux I__8041 (
            .O(N__39932),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ));
    InMux I__8040 (
            .O(N__39927),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ));
    InMux I__8039 (
            .O(N__39924),
            .I(N__39920));
    InMux I__8038 (
            .O(N__39923),
            .I(N__39917));
    LocalMux I__8037 (
            .O(N__39920),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ));
    LocalMux I__8036 (
            .O(N__39917),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ));
    InMux I__8035 (
            .O(N__39912),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ));
    InMux I__8034 (
            .O(N__39909),
            .I(N__39903));
    InMux I__8033 (
            .O(N__39908),
            .I(N__39903));
    LocalMux I__8032 (
            .O(N__39903),
            .I(N__39899));
    InMux I__8031 (
            .O(N__39902),
            .I(N__39896));
    Span4Mux_v I__8030 (
            .O(N__39899),
            .I(N__39893));
    LocalMux I__8029 (
            .O(N__39896),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ));
    Odrv4 I__8028 (
            .O(N__39893),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ));
    InMux I__8027 (
            .O(N__39888),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_27 ));
    CascadeMux I__8026 (
            .O(N__39885),
            .I(N__39882));
    InMux I__8025 (
            .O(N__39882),
            .I(N__39876));
    InMux I__8024 (
            .O(N__39881),
            .I(N__39876));
    LocalMux I__8023 (
            .O(N__39876),
            .I(N__39872));
    InMux I__8022 (
            .O(N__39875),
            .I(N__39869));
    Span4Mux_v I__8021 (
            .O(N__39872),
            .I(N__39866));
    LocalMux I__8020 (
            .O(N__39869),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ));
    Odrv4 I__8019 (
            .O(N__39866),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ));
    InMux I__8018 (
            .O(N__39861),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_28 ));
    InMux I__8017 (
            .O(N__39858),
            .I(N__39854));
    InMux I__8016 (
            .O(N__39857),
            .I(N__39851));
    LocalMux I__8015 (
            .O(N__39854),
            .I(N__39845));
    LocalMux I__8014 (
            .O(N__39851),
            .I(N__39845));
    InMux I__8013 (
            .O(N__39850),
            .I(N__39842));
    Span4Mux_v I__8012 (
            .O(N__39845),
            .I(N__39839));
    LocalMux I__8011 (
            .O(N__39842),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    Odrv4 I__8010 (
            .O(N__39839),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    InMux I__8009 (
            .O(N__39834),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_29 ));
    InMux I__8008 (
            .O(N__39831),
            .I(N__39791));
    InMux I__8007 (
            .O(N__39830),
            .I(N__39791));
    InMux I__8006 (
            .O(N__39829),
            .I(N__39791));
    InMux I__8005 (
            .O(N__39828),
            .I(N__39791));
    InMux I__8004 (
            .O(N__39827),
            .I(N__39782));
    InMux I__8003 (
            .O(N__39826),
            .I(N__39782));
    InMux I__8002 (
            .O(N__39825),
            .I(N__39782));
    InMux I__8001 (
            .O(N__39824),
            .I(N__39782));
    InMux I__8000 (
            .O(N__39823),
            .I(N__39773));
    InMux I__7999 (
            .O(N__39822),
            .I(N__39773));
    InMux I__7998 (
            .O(N__39821),
            .I(N__39773));
    InMux I__7997 (
            .O(N__39820),
            .I(N__39773));
    InMux I__7996 (
            .O(N__39819),
            .I(N__39764));
    InMux I__7995 (
            .O(N__39818),
            .I(N__39764));
    InMux I__7994 (
            .O(N__39817),
            .I(N__39764));
    InMux I__7993 (
            .O(N__39816),
            .I(N__39764));
    InMux I__7992 (
            .O(N__39815),
            .I(N__39755));
    InMux I__7991 (
            .O(N__39814),
            .I(N__39755));
    InMux I__7990 (
            .O(N__39813),
            .I(N__39755));
    InMux I__7989 (
            .O(N__39812),
            .I(N__39755));
    InMux I__7988 (
            .O(N__39811),
            .I(N__39746));
    InMux I__7987 (
            .O(N__39810),
            .I(N__39746));
    InMux I__7986 (
            .O(N__39809),
            .I(N__39746));
    InMux I__7985 (
            .O(N__39808),
            .I(N__39746));
    InMux I__7984 (
            .O(N__39807),
            .I(N__39737));
    InMux I__7983 (
            .O(N__39806),
            .I(N__39737));
    InMux I__7982 (
            .O(N__39805),
            .I(N__39737));
    InMux I__7981 (
            .O(N__39804),
            .I(N__39737));
    InMux I__7980 (
            .O(N__39803),
            .I(N__39728));
    InMux I__7979 (
            .O(N__39802),
            .I(N__39728));
    InMux I__7978 (
            .O(N__39801),
            .I(N__39728));
    InMux I__7977 (
            .O(N__39800),
            .I(N__39728));
    LocalMux I__7976 (
            .O(N__39791),
            .I(N__39723));
    LocalMux I__7975 (
            .O(N__39782),
            .I(N__39723));
    LocalMux I__7974 (
            .O(N__39773),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    LocalMux I__7973 (
            .O(N__39764),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    LocalMux I__7972 (
            .O(N__39755),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    LocalMux I__7971 (
            .O(N__39746),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    LocalMux I__7970 (
            .O(N__39737),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    LocalMux I__7969 (
            .O(N__39728),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    Odrv4 I__7968 (
            .O(N__39723),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    InMux I__7967 (
            .O(N__39708),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_30 ));
    InMux I__7966 (
            .O(N__39705),
            .I(N__39701));
    InMux I__7965 (
            .O(N__39704),
            .I(N__39698));
    LocalMux I__7964 (
            .O(N__39701),
            .I(N__39692));
    LocalMux I__7963 (
            .O(N__39698),
            .I(N__39692));
    InMux I__7962 (
            .O(N__39697),
            .I(N__39689));
    Span4Mux_v I__7961 (
            .O(N__39692),
            .I(N__39686));
    LocalMux I__7960 (
            .O(N__39689),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    Odrv4 I__7959 (
            .O(N__39686),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    CEMux I__7958 (
            .O(N__39681),
            .I(N__39676));
    CEMux I__7957 (
            .O(N__39680),
            .I(N__39672));
    CEMux I__7956 (
            .O(N__39679),
            .I(N__39669));
    LocalMux I__7955 (
            .O(N__39676),
            .I(N__39666));
    CEMux I__7954 (
            .O(N__39675),
            .I(N__39663));
    LocalMux I__7953 (
            .O(N__39672),
            .I(N__39660));
    LocalMux I__7952 (
            .O(N__39669),
            .I(N__39657));
    Span4Mux_v I__7951 (
            .O(N__39666),
            .I(N__39654));
    LocalMux I__7950 (
            .O(N__39663),
            .I(N__39649));
    Span4Mux_v I__7949 (
            .O(N__39660),
            .I(N__39649));
    Span4Mux_v I__7948 (
            .O(N__39657),
            .I(N__39646));
    Span4Mux_h I__7947 (
            .O(N__39654),
            .I(N__39641));
    Span4Mux_v I__7946 (
            .O(N__39649),
            .I(N__39641));
    Span4Mux_h I__7945 (
            .O(N__39646),
            .I(N__39638));
    Span4Mux_h I__7944 (
            .O(N__39641),
            .I(N__39635));
    Odrv4 I__7943 (
            .O(N__39638),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__7942 (
            .O(N__39635),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__7941 (
            .O(N__39630),
            .I(N__39627));
    InMux I__7940 (
            .O(N__39627),
            .I(N__39624));
    LocalMux I__7939 (
            .O(N__39624),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ));
    InMux I__7938 (
            .O(N__39621),
            .I(N__39618));
    LocalMux I__7937 (
            .O(N__39618),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ));
    InMux I__7936 (
            .O(N__39615),
            .I(N__39611));
    InMux I__7935 (
            .O(N__39614),
            .I(N__39608));
    LocalMux I__7934 (
            .O(N__39611),
            .I(N__39605));
    LocalMux I__7933 (
            .O(N__39608),
            .I(N__39601));
    Span4Mux_v I__7932 (
            .O(N__39605),
            .I(N__39598));
    CascadeMux I__7931 (
            .O(N__39604),
            .I(N__39595));
    Span4Mux_v I__7930 (
            .O(N__39601),
            .I(N__39590));
    Span4Mux_v I__7929 (
            .O(N__39598),
            .I(N__39590));
    InMux I__7928 (
            .O(N__39595),
            .I(N__39587));
    Odrv4 I__7927 (
            .O(N__39590),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ));
    LocalMux I__7926 (
            .O(N__39587),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ));
    InMux I__7925 (
            .O(N__39582),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ));
    InMux I__7924 (
            .O(N__39579),
            .I(N__39575));
    InMux I__7923 (
            .O(N__39578),
            .I(N__39572));
    LocalMux I__7922 (
            .O(N__39575),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ));
    LocalMux I__7921 (
            .O(N__39572),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ));
    InMux I__7920 (
            .O(N__39567),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ));
    InMux I__7919 (
            .O(N__39564),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_18 ));
    InMux I__7918 (
            .O(N__39561),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_19 ));
    InMux I__7917 (
            .O(N__39558),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_20 ));
    InMux I__7916 (
            .O(N__39555),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_21 ));
    InMux I__7915 (
            .O(N__39552),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_22 ));
    InMux I__7914 (
            .O(N__39549),
            .I(bfn_14_19_0_));
    InMux I__7913 (
            .O(N__39546),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_24 ));
    InMux I__7912 (
            .O(N__39543),
            .I(N__39536));
    InMux I__7911 (
            .O(N__39542),
            .I(N__39536));
    InMux I__7910 (
            .O(N__39541),
            .I(N__39533));
    LocalMux I__7909 (
            .O(N__39536),
            .I(N__39530));
    LocalMux I__7908 (
            .O(N__39533),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ));
    Odrv12 I__7907 (
            .O(N__39530),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ));
    InMux I__7906 (
            .O(N__39525),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_25 ));
    InMux I__7905 (
            .O(N__39522),
            .I(N__39516));
    InMux I__7904 (
            .O(N__39521),
            .I(N__39516));
    LocalMux I__7903 (
            .O(N__39516),
            .I(N__39512));
    InMux I__7902 (
            .O(N__39515),
            .I(N__39509));
    Span4Mux_h I__7901 (
            .O(N__39512),
            .I(N__39506));
    LocalMux I__7900 (
            .O(N__39509),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ));
    Odrv4 I__7899 (
            .O(N__39506),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ));
    InMux I__7898 (
            .O(N__39501),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_26 ));
    InMux I__7897 (
            .O(N__39498),
            .I(N__39494));
    InMux I__7896 (
            .O(N__39497),
            .I(N__39491));
    LocalMux I__7895 (
            .O(N__39494),
            .I(N__39488));
    LocalMux I__7894 (
            .O(N__39491),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ));
    Odrv12 I__7893 (
            .O(N__39488),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ));
    InMux I__7892 (
            .O(N__39483),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_9 ));
    InMux I__7891 (
            .O(N__39480),
            .I(N__39476));
    InMux I__7890 (
            .O(N__39479),
            .I(N__39473));
    LocalMux I__7889 (
            .O(N__39476),
            .I(N__39470));
    LocalMux I__7888 (
            .O(N__39473),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ));
    Odrv12 I__7887 (
            .O(N__39470),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ));
    InMux I__7886 (
            .O(N__39465),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_10 ));
    InMux I__7885 (
            .O(N__39462),
            .I(N__39459));
    LocalMux I__7884 (
            .O(N__39459),
            .I(N__39455));
    InMux I__7883 (
            .O(N__39458),
            .I(N__39452));
    Span4Mux_v I__7882 (
            .O(N__39455),
            .I(N__39449));
    LocalMux I__7881 (
            .O(N__39452),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ));
    Odrv4 I__7880 (
            .O(N__39449),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ));
    InMux I__7879 (
            .O(N__39444),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_11 ));
    InMux I__7878 (
            .O(N__39441),
            .I(N__39437));
    InMux I__7877 (
            .O(N__39440),
            .I(N__39434));
    LocalMux I__7876 (
            .O(N__39437),
            .I(N__39431));
    LocalMux I__7875 (
            .O(N__39434),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ));
    Odrv12 I__7874 (
            .O(N__39431),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ));
    InMux I__7873 (
            .O(N__39426),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_12 ));
    InMux I__7872 (
            .O(N__39423),
            .I(N__39419));
    InMux I__7871 (
            .O(N__39422),
            .I(N__39416));
    LocalMux I__7870 (
            .O(N__39419),
            .I(N__39413));
    LocalMux I__7869 (
            .O(N__39416),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ));
    Odrv12 I__7868 (
            .O(N__39413),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ));
    InMux I__7867 (
            .O(N__39408),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_13 ));
    InMux I__7866 (
            .O(N__39405),
            .I(N__39401));
    InMux I__7865 (
            .O(N__39404),
            .I(N__39398));
    LocalMux I__7864 (
            .O(N__39401),
            .I(N__39395));
    LocalMux I__7863 (
            .O(N__39398),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ));
    Odrv12 I__7862 (
            .O(N__39395),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ));
    InMux I__7861 (
            .O(N__39390),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_14 ));
    InMux I__7860 (
            .O(N__39387),
            .I(bfn_14_18_0_));
    InMux I__7859 (
            .O(N__39384),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_16 ));
    InMux I__7858 (
            .O(N__39381),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_17 ));
    InMux I__7857 (
            .O(N__39378),
            .I(N__39374));
    InMux I__7856 (
            .O(N__39377),
            .I(N__39371));
    LocalMux I__7855 (
            .O(N__39374),
            .I(N__39368));
    LocalMux I__7854 (
            .O(N__39371),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ));
    Odrv12 I__7853 (
            .O(N__39368),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ));
    InMux I__7852 (
            .O(N__39363),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_1 ));
    InMux I__7851 (
            .O(N__39360),
            .I(N__39356));
    InMux I__7850 (
            .O(N__39359),
            .I(N__39353));
    LocalMux I__7849 (
            .O(N__39356),
            .I(N__39350));
    LocalMux I__7848 (
            .O(N__39353),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ));
    Odrv12 I__7847 (
            .O(N__39350),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ));
    InMux I__7846 (
            .O(N__39345),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_2 ));
    InMux I__7845 (
            .O(N__39342),
            .I(N__39338));
    InMux I__7844 (
            .O(N__39341),
            .I(N__39335));
    LocalMux I__7843 (
            .O(N__39338),
            .I(N__39332));
    LocalMux I__7842 (
            .O(N__39335),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ));
    Odrv12 I__7841 (
            .O(N__39332),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ));
    InMux I__7840 (
            .O(N__39327),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_3 ));
    InMux I__7839 (
            .O(N__39324),
            .I(N__39320));
    InMux I__7838 (
            .O(N__39323),
            .I(N__39317));
    LocalMux I__7837 (
            .O(N__39320),
            .I(N__39314));
    LocalMux I__7836 (
            .O(N__39317),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ));
    Odrv12 I__7835 (
            .O(N__39314),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ));
    InMux I__7834 (
            .O(N__39309),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_4 ));
    InMux I__7833 (
            .O(N__39306),
            .I(N__39302));
    InMux I__7832 (
            .O(N__39305),
            .I(N__39299));
    LocalMux I__7831 (
            .O(N__39302),
            .I(N__39296));
    LocalMux I__7830 (
            .O(N__39299),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ));
    Odrv12 I__7829 (
            .O(N__39296),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ));
    InMux I__7828 (
            .O(N__39291),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_5 ));
    InMux I__7827 (
            .O(N__39288),
            .I(N__39284));
    InMux I__7826 (
            .O(N__39287),
            .I(N__39281));
    LocalMux I__7825 (
            .O(N__39284),
            .I(N__39278));
    LocalMux I__7824 (
            .O(N__39281),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ));
    Odrv12 I__7823 (
            .O(N__39278),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ));
    InMux I__7822 (
            .O(N__39273),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_6 ));
    InMux I__7821 (
            .O(N__39270),
            .I(N__39266));
    InMux I__7820 (
            .O(N__39269),
            .I(N__39263));
    LocalMux I__7819 (
            .O(N__39266),
            .I(N__39260));
    LocalMux I__7818 (
            .O(N__39263),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ));
    Odrv12 I__7817 (
            .O(N__39260),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ));
    InMux I__7816 (
            .O(N__39255),
            .I(bfn_14_17_0_));
    InMux I__7815 (
            .O(N__39252),
            .I(N__39248));
    InMux I__7814 (
            .O(N__39251),
            .I(N__39245));
    LocalMux I__7813 (
            .O(N__39248),
            .I(N__39242));
    LocalMux I__7812 (
            .O(N__39245),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ));
    Odrv12 I__7811 (
            .O(N__39242),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ));
    InMux I__7810 (
            .O(N__39237),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_8 ));
    InMux I__7809 (
            .O(N__39234),
            .I(bfn_14_15_0_));
    CascadeMux I__7808 (
            .O(N__39231),
            .I(N__39227));
    InMux I__7807 (
            .O(N__39230),
            .I(N__39222));
    InMux I__7806 (
            .O(N__39227),
            .I(N__39222));
    LocalMux I__7805 (
            .O(N__39222),
            .I(N__39219));
    Span4Mux_h I__7804 (
            .O(N__39219),
            .I(N__39216));
    Odrv4 I__7803 (
            .O(N__39216),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ));
    CascadeMux I__7802 (
            .O(N__39213),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO_cascade_ ));
    InMux I__7801 (
            .O(N__39210),
            .I(N__39204));
    InMux I__7800 (
            .O(N__39209),
            .I(N__39201));
    InMux I__7799 (
            .O(N__39208),
            .I(N__39198));
    CascadeMux I__7798 (
            .O(N__39207),
            .I(N__39194));
    LocalMux I__7797 (
            .O(N__39204),
            .I(N__39190));
    LocalMux I__7796 (
            .O(N__39201),
            .I(N__39187));
    LocalMux I__7795 (
            .O(N__39198),
            .I(N__39184));
    InMux I__7794 (
            .O(N__39197),
            .I(N__39181));
    InMux I__7793 (
            .O(N__39194),
            .I(N__39176));
    InMux I__7792 (
            .O(N__39193),
            .I(N__39176));
    Span4Mux_v I__7791 (
            .O(N__39190),
            .I(N__39173));
    Span4Mux_v I__7790 (
            .O(N__39187),
            .I(N__39168));
    Span4Mux_v I__7789 (
            .O(N__39184),
            .I(N__39168));
    LocalMux I__7788 (
            .O(N__39181),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__7787 (
            .O(N__39176),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7786 (
            .O(N__39173),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7785 (
            .O(N__39168),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__7784 (
            .O(N__39159),
            .I(N__39153));
    InMux I__7783 (
            .O(N__39158),
            .I(N__39150));
    InMux I__7782 (
            .O(N__39157),
            .I(N__39145));
    InMux I__7781 (
            .O(N__39156),
            .I(N__39145));
    LocalMux I__7780 (
            .O(N__39153),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ));
    LocalMux I__7779 (
            .O(N__39150),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ));
    LocalMux I__7778 (
            .O(N__39145),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ));
    CascadeMux I__7777 (
            .O(N__39138),
            .I(N__39135));
    InMux I__7776 (
            .O(N__39135),
            .I(N__39132));
    LocalMux I__7775 (
            .O(N__39132),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt30 ));
    CascadeMux I__7774 (
            .O(N__39129),
            .I(N__39126));
    InMux I__7773 (
            .O(N__39126),
            .I(N__39123));
    LocalMux I__7772 (
            .O(N__39123),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt26 ));
    InMux I__7771 (
            .O(N__39120),
            .I(N__39117));
    LocalMux I__7770 (
            .O(N__39117),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ));
    InMux I__7769 (
            .O(N__39114),
            .I(N__39111));
    LocalMux I__7768 (
            .O(N__39111),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    CascadeMux I__7767 (
            .O(N__39108),
            .I(elapsed_time_ns_1_RNILK91B_0_9_cascade_));
    InMux I__7766 (
            .O(N__39105),
            .I(N__39101));
    CascadeMux I__7765 (
            .O(N__39104),
            .I(N__39098));
    LocalMux I__7764 (
            .O(N__39101),
            .I(N__39095));
    InMux I__7763 (
            .O(N__39098),
            .I(N__39092));
    Odrv4 I__7762 (
            .O(N__39095),
            .I(\phase_controller_inst1.stoper_hc.counter ));
    LocalMux I__7761 (
            .O(N__39092),
            .I(\phase_controller_inst1.stoper_hc.counter ));
    InMux I__7760 (
            .O(N__39087),
            .I(N__39083));
    InMux I__7759 (
            .O(N__39086),
            .I(N__39080));
    LocalMux I__7758 (
            .O(N__39083),
            .I(N__39077));
    LocalMux I__7757 (
            .O(N__39080),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ));
    Odrv12 I__7756 (
            .O(N__39077),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ));
    InMux I__7755 (
            .O(N__39072),
            .I(N__39068));
    InMux I__7754 (
            .O(N__39071),
            .I(N__39065));
    LocalMux I__7753 (
            .O(N__39068),
            .I(N__39062));
    LocalMux I__7752 (
            .O(N__39065),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ));
    Odrv12 I__7751 (
            .O(N__39062),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ));
    InMux I__7750 (
            .O(N__39057),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_0 ));
    CascadeMux I__7749 (
            .O(N__39054),
            .I(N__39051));
    InMux I__7748 (
            .O(N__39051),
            .I(N__39048));
    LocalMux I__7747 (
            .O(N__39048),
            .I(\phase_controller_inst1.stoper_hc.counter_i_15 ));
    InMux I__7746 (
            .O(N__39045),
            .I(N__39042));
    LocalMux I__7745 (
            .O(N__39042),
            .I(N__39039));
    Odrv4 I__7744 (
            .O(N__39039),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ));
    InMux I__7743 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__7742 (
            .O(N__39033),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ));
    CascadeMux I__7741 (
            .O(N__39030),
            .I(N__39027));
    InMux I__7740 (
            .O(N__39027),
            .I(N__39024));
    LocalMux I__7739 (
            .O(N__39024),
            .I(N__39021));
    Odrv4 I__7738 (
            .O(N__39021),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt28 ));
    InMux I__7737 (
            .O(N__39018),
            .I(N__39015));
    LocalMux I__7736 (
            .O(N__39015),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__7735 (
            .O(N__39012),
            .I(N__39009));
    InMux I__7734 (
            .O(N__39009),
            .I(N__39006));
    LocalMux I__7733 (
            .O(N__39006),
            .I(\phase_controller_inst1.stoper_hc.counter_i_7 ));
    CascadeMux I__7732 (
            .O(N__39003),
            .I(N__39000));
    InMux I__7731 (
            .O(N__39000),
            .I(N__38997));
    LocalMux I__7730 (
            .O(N__38997),
            .I(\phase_controller_inst1.stoper_hc.counter_i_8 ));
    CascadeMux I__7729 (
            .O(N__38994),
            .I(N__38991));
    InMux I__7728 (
            .O(N__38991),
            .I(N__38988));
    LocalMux I__7727 (
            .O(N__38988),
            .I(\phase_controller_inst1.stoper_hc.counter_i_9 ));
    CascadeMux I__7726 (
            .O(N__38985),
            .I(N__38982));
    InMux I__7725 (
            .O(N__38982),
            .I(N__38979));
    LocalMux I__7724 (
            .O(N__38979),
            .I(\phase_controller_inst1.stoper_hc.counter_i_10 ));
    CascadeMux I__7723 (
            .O(N__38976),
            .I(N__38973));
    InMux I__7722 (
            .O(N__38973),
            .I(N__38970));
    LocalMux I__7721 (
            .O(N__38970),
            .I(N__38967));
    Odrv4 I__7720 (
            .O(N__38967),
            .I(\phase_controller_inst1.stoper_hc.counter_i_11 ));
    CascadeMux I__7719 (
            .O(N__38964),
            .I(N__38961));
    InMux I__7718 (
            .O(N__38961),
            .I(N__38958));
    LocalMux I__7717 (
            .O(N__38958),
            .I(N__38955));
    Odrv4 I__7716 (
            .O(N__38955),
            .I(\phase_controller_inst1.stoper_hc.counter_i_12 ));
    CascadeMux I__7715 (
            .O(N__38952),
            .I(N__38949));
    InMux I__7714 (
            .O(N__38949),
            .I(N__38946));
    LocalMux I__7713 (
            .O(N__38946),
            .I(\phase_controller_inst1.stoper_hc.counter_i_13 ));
    CascadeMux I__7712 (
            .O(N__38943),
            .I(N__38940));
    InMux I__7711 (
            .O(N__38940),
            .I(N__38937));
    LocalMux I__7710 (
            .O(N__38937),
            .I(\phase_controller_inst1.stoper_hc.counter_i_14 ));
    InMux I__7709 (
            .O(N__38934),
            .I(N__38929));
    InMux I__7708 (
            .O(N__38933),
            .I(N__38924));
    InMux I__7707 (
            .O(N__38932),
            .I(N__38924));
    LocalMux I__7706 (
            .O(N__38929),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ));
    LocalMux I__7705 (
            .O(N__38924),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ));
    CascadeMux I__7704 (
            .O(N__38919),
            .I(N__38915));
    InMux I__7703 (
            .O(N__38918),
            .I(N__38908));
    InMux I__7702 (
            .O(N__38915),
            .I(N__38908));
    InMux I__7701 (
            .O(N__38914),
            .I(N__38903));
    InMux I__7700 (
            .O(N__38913),
            .I(N__38903));
    LocalMux I__7699 (
            .O(N__38908),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ));
    LocalMux I__7698 (
            .O(N__38903),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ));
    InMux I__7697 (
            .O(N__38898),
            .I(N__38893));
    InMux I__7696 (
            .O(N__38897),
            .I(N__38888));
    InMux I__7695 (
            .O(N__38896),
            .I(N__38888));
    LocalMux I__7694 (
            .O(N__38893),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ));
    LocalMux I__7693 (
            .O(N__38888),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ));
    InMux I__7692 (
            .O(N__38883),
            .I(N__38880));
    LocalMux I__7691 (
            .O(N__38880),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt28 ));
    InMux I__7690 (
            .O(N__38877),
            .I(N__38874));
    LocalMux I__7689 (
            .O(N__38874),
            .I(N__38871));
    Span4Mux_v I__7688 (
            .O(N__38871),
            .I(N__38868));
    Span4Mux_h I__7687 (
            .O(N__38868),
            .I(N__38865));
    Odrv4 I__7686 (
            .O(N__38865),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ));
    CascadeMux I__7685 (
            .O(N__38862),
            .I(N__38859));
    InMux I__7684 (
            .O(N__38859),
            .I(N__38856));
    LocalMux I__7683 (
            .O(N__38856),
            .I(\phase_controller_inst1.stoper_hc.counter_i_0 ));
    CascadeMux I__7682 (
            .O(N__38853),
            .I(N__38850));
    InMux I__7681 (
            .O(N__38850),
            .I(N__38847));
    LocalMux I__7680 (
            .O(N__38847),
            .I(\phase_controller_inst1.stoper_hc.counter_i_1 ));
    CascadeMux I__7679 (
            .O(N__38844),
            .I(N__38841));
    InMux I__7678 (
            .O(N__38841),
            .I(N__38838));
    LocalMux I__7677 (
            .O(N__38838),
            .I(\phase_controller_inst1.stoper_hc.counter_i_2 ));
    CascadeMux I__7676 (
            .O(N__38835),
            .I(N__38832));
    InMux I__7675 (
            .O(N__38832),
            .I(N__38829));
    LocalMux I__7674 (
            .O(N__38829),
            .I(\phase_controller_inst1.stoper_hc.counter_i_3 ));
    CascadeMux I__7673 (
            .O(N__38826),
            .I(N__38823));
    InMux I__7672 (
            .O(N__38823),
            .I(N__38820));
    LocalMux I__7671 (
            .O(N__38820),
            .I(N__38817));
    Odrv4 I__7670 (
            .O(N__38817),
            .I(\phase_controller_inst1.stoper_hc.counter_i_4 ));
    CascadeMux I__7669 (
            .O(N__38814),
            .I(N__38811));
    InMux I__7668 (
            .O(N__38811),
            .I(N__38808));
    LocalMux I__7667 (
            .O(N__38808),
            .I(\phase_controller_inst1.stoper_hc.counter_i_5 ));
    CascadeMux I__7666 (
            .O(N__38805),
            .I(N__38802));
    InMux I__7665 (
            .O(N__38802),
            .I(N__38799));
    LocalMux I__7664 (
            .O(N__38799),
            .I(\phase_controller_inst1.stoper_hc.counter_i_6 ));
    InMux I__7663 (
            .O(N__38796),
            .I(N__38793));
    LocalMux I__7662 (
            .O(N__38793),
            .I(N__38790));
    Odrv4 I__7661 (
            .O(N__38790),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ));
    CascadeMux I__7660 (
            .O(N__38787),
            .I(N__38784));
    InMux I__7659 (
            .O(N__38784),
            .I(N__38781));
    LocalMux I__7658 (
            .O(N__38781),
            .I(N__38778));
    Odrv4 I__7657 (
            .O(N__38778),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt30 ));
    InMux I__7656 (
            .O(N__38775),
            .I(bfn_14_11_0_));
    InMux I__7655 (
            .O(N__38772),
            .I(N__38766));
    InMux I__7654 (
            .O(N__38771),
            .I(N__38766));
    LocalMux I__7653 (
            .O(N__38766),
            .I(N__38763));
    Span4Mux_v I__7652 (
            .O(N__38763),
            .I(N__38759));
    InMux I__7651 (
            .O(N__38762),
            .I(N__38756));
    Span4Mux_h I__7650 (
            .O(N__38759),
            .I(N__38753));
    LocalMux I__7649 (
            .O(N__38756),
            .I(N__38750));
    Odrv4 I__7648 (
            .O(N__38753),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    Odrv12 I__7647 (
            .O(N__38750),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    CascadeMux I__7646 (
            .O(N__38745),
            .I(N__38742));
    InMux I__7645 (
            .O(N__38742),
            .I(N__38739));
    LocalMux I__7644 (
            .O(N__38739),
            .I(N__38736));
    Odrv4 I__7643 (
            .O(N__38736),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ));
    InMux I__7642 (
            .O(N__38733),
            .I(N__38729));
    InMux I__7641 (
            .O(N__38732),
            .I(N__38726));
    LocalMux I__7640 (
            .O(N__38729),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ));
    LocalMux I__7639 (
            .O(N__38726),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ));
    CascadeMux I__7638 (
            .O(N__38721),
            .I(N__38718));
    InMux I__7637 (
            .O(N__38718),
            .I(N__38715));
    LocalMux I__7636 (
            .O(N__38715),
            .I(\phase_controller_inst2.stoper_hc.counter_i_10 ));
    InMux I__7635 (
            .O(N__38712),
            .I(N__38708));
    InMux I__7634 (
            .O(N__38711),
            .I(N__38705));
    LocalMux I__7633 (
            .O(N__38708),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ));
    LocalMux I__7632 (
            .O(N__38705),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ));
    CascadeMux I__7631 (
            .O(N__38700),
            .I(N__38697));
    InMux I__7630 (
            .O(N__38697),
            .I(N__38694));
    LocalMux I__7629 (
            .O(N__38694),
            .I(\phase_controller_inst2.stoper_hc.counter_i_11 ));
    InMux I__7628 (
            .O(N__38691),
            .I(N__38687));
    InMux I__7627 (
            .O(N__38690),
            .I(N__38684));
    LocalMux I__7626 (
            .O(N__38687),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ));
    LocalMux I__7625 (
            .O(N__38684),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ));
    CascadeMux I__7624 (
            .O(N__38679),
            .I(N__38676));
    InMux I__7623 (
            .O(N__38676),
            .I(N__38673));
    LocalMux I__7622 (
            .O(N__38673),
            .I(N__38670));
    Odrv4 I__7621 (
            .O(N__38670),
            .I(\phase_controller_inst2.stoper_hc.counter_i_12 ));
    InMux I__7620 (
            .O(N__38667),
            .I(N__38663));
    InMux I__7619 (
            .O(N__38666),
            .I(N__38660));
    LocalMux I__7618 (
            .O(N__38663),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ));
    LocalMux I__7617 (
            .O(N__38660),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ));
    CascadeMux I__7616 (
            .O(N__38655),
            .I(N__38652));
    InMux I__7615 (
            .O(N__38652),
            .I(N__38649));
    LocalMux I__7614 (
            .O(N__38649),
            .I(\phase_controller_inst2.stoper_hc.counter_i_13 ));
    InMux I__7613 (
            .O(N__38646),
            .I(N__38642));
    InMux I__7612 (
            .O(N__38645),
            .I(N__38639));
    LocalMux I__7611 (
            .O(N__38642),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ));
    LocalMux I__7610 (
            .O(N__38639),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ));
    CascadeMux I__7609 (
            .O(N__38634),
            .I(N__38631));
    InMux I__7608 (
            .O(N__38631),
            .I(N__38628));
    LocalMux I__7607 (
            .O(N__38628),
            .I(\phase_controller_inst2.stoper_hc.counter_i_14 ));
    InMux I__7606 (
            .O(N__38625),
            .I(N__38621));
    InMux I__7605 (
            .O(N__38624),
            .I(N__38618));
    LocalMux I__7604 (
            .O(N__38621),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ));
    LocalMux I__7603 (
            .O(N__38618),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ));
    CascadeMux I__7602 (
            .O(N__38613),
            .I(N__38610));
    InMux I__7601 (
            .O(N__38610),
            .I(N__38607));
    LocalMux I__7600 (
            .O(N__38607),
            .I(\phase_controller_inst2.stoper_hc.counter_i_15 ));
    InMux I__7599 (
            .O(N__38604),
            .I(N__38600));
    InMux I__7598 (
            .O(N__38603),
            .I(N__38597));
    LocalMux I__7597 (
            .O(N__38600),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ));
    LocalMux I__7596 (
            .O(N__38597),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ));
    InMux I__7595 (
            .O(N__38592),
            .I(N__38589));
    LocalMux I__7594 (
            .O(N__38589),
            .I(\phase_controller_inst2.stoper_hc.counter_i_2 ));
    InMux I__7593 (
            .O(N__38586),
            .I(N__38582));
    InMux I__7592 (
            .O(N__38585),
            .I(N__38579));
    LocalMux I__7591 (
            .O(N__38582),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ));
    LocalMux I__7590 (
            .O(N__38579),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ));
    InMux I__7589 (
            .O(N__38574),
            .I(N__38571));
    LocalMux I__7588 (
            .O(N__38571),
            .I(\phase_controller_inst2.stoper_hc.counter_i_3 ));
    InMux I__7587 (
            .O(N__38568),
            .I(N__38564));
    InMux I__7586 (
            .O(N__38567),
            .I(N__38561));
    LocalMux I__7585 (
            .O(N__38564),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ));
    LocalMux I__7584 (
            .O(N__38561),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ));
    InMux I__7583 (
            .O(N__38556),
            .I(N__38553));
    LocalMux I__7582 (
            .O(N__38553),
            .I(\phase_controller_inst2.stoper_hc.counter_i_4 ));
    InMux I__7581 (
            .O(N__38550),
            .I(N__38546));
    InMux I__7580 (
            .O(N__38549),
            .I(N__38543));
    LocalMux I__7579 (
            .O(N__38546),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ));
    LocalMux I__7578 (
            .O(N__38543),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ));
    CascadeMux I__7577 (
            .O(N__38538),
            .I(N__38535));
    InMux I__7576 (
            .O(N__38535),
            .I(N__38532));
    LocalMux I__7575 (
            .O(N__38532),
            .I(\phase_controller_inst2.stoper_hc.counter_i_5 ));
    InMux I__7574 (
            .O(N__38529),
            .I(N__38525));
    InMux I__7573 (
            .O(N__38528),
            .I(N__38522));
    LocalMux I__7572 (
            .O(N__38525),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ));
    LocalMux I__7571 (
            .O(N__38522),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ));
    CascadeMux I__7570 (
            .O(N__38517),
            .I(N__38514));
    InMux I__7569 (
            .O(N__38514),
            .I(N__38511));
    LocalMux I__7568 (
            .O(N__38511),
            .I(N__38508));
    Odrv4 I__7567 (
            .O(N__38508),
            .I(\phase_controller_inst2.stoper_hc.counter_i_6 ));
    InMux I__7566 (
            .O(N__38505),
            .I(N__38501));
    InMux I__7565 (
            .O(N__38504),
            .I(N__38498));
    LocalMux I__7564 (
            .O(N__38501),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ));
    LocalMux I__7563 (
            .O(N__38498),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ));
    CascadeMux I__7562 (
            .O(N__38493),
            .I(N__38490));
    InMux I__7561 (
            .O(N__38490),
            .I(N__38487));
    LocalMux I__7560 (
            .O(N__38487),
            .I(\phase_controller_inst2.stoper_hc.counter_i_7 ));
    InMux I__7559 (
            .O(N__38484),
            .I(N__38480));
    InMux I__7558 (
            .O(N__38483),
            .I(N__38477));
    LocalMux I__7557 (
            .O(N__38480),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ));
    LocalMux I__7556 (
            .O(N__38477),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ));
    CascadeMux I__7555 (
            .O(N__38472),
            .I(N__38469));
    InMux I__7554 (
            .O(N__38469),
            .I(N__38466));
    LocalMux I__7553 (
            .O(N__38466),
            .I(\phase_controller_inst2.stoper_hc.counter_i_8 ));
    InMux I__7552 (
            .O(N__38463),
            .I(N__38459));
    InMux I__7551 (
            .O(N__38462),
            .I(N__38456));
    LocalMux I__7550 (
            .O(N__38459),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ));
    LocalMux I__7549 (
            .O(N__38456),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ));
    CascadeMux I__7548 (
            .O(N__38451),
            .I(N__38448));
    InMux I__7547 (
            .O(N__38448),
            .I(N__38445));
    LocalMux I__7546 (
            .O(N__38445),
            .I(\phase_controller_inst2.stoper_hc.counter_i_9 ));
    InMux I__7545 (
            .O(N__38442),
            .I(N__38438));
    InMux I__7544 (
            .O(N__38441),
            .I(N__38435));
    LocalMux I__7543 (
            .O(N__38438),
            .I(N__38432));
    LocalMux I__7542 (
            .O(N__38435),
            .I(N__38429));
    Odrv12 I__7541 (
            .O(N__38432),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_19));
    Odrv12 I__7540 (
            .O(N__38429),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_19));
    CEMux I__7539 (
            .O(N__38424),
            .I(N__38420));
    CEMux I__7538 (
            .O(N__38423),
            .I(N__38416));
    LocalMux I__7537 (
            .O(N__38420),
            .I(N__38413));
    CEMux I__7536 (
            .O(N__38419),
            .I(N__38410));
    LocalMux I__7535 (
            .O(N__38416),
            .I(N__38406));
    Span4Mux_h I__7534 (
            .O(N__38413),
            .I(N__38401));
    LocalMux I__7533 (
            .O(N__38410),
            .I(N__38398));
    CEMux I__7532 (
            .O(N__38409),
            .I(N__38395));
    Span4Mux_v I__7531 (
            .O(N__38406),
            .I(N__38392));
    CEMux I__7530 (
            .O(N__38405),
            .I(N__38389));
    CEMux I__7529 (
            .O(N__38404),
            .I(N__38386));
    Span4Mux_v I__7528 (
            .O(N__38401),
            .I(N__38375));
    Span4Mux_v I__7527 (
            .O(N__38398),
            .I(N__38375));
    LocalMux I__7526 (
            .O(N__38395),
            .I(N__38375));
    Span4Mux_v I__7525 (
            .O(N__38392),
            .I(N__38375));
    LocalMux I__7524 (
            .O(N__38389),
            .I(N__38375));
    LocalMux I__7523 (
            .O(N__38386),
            .I(N__38371));
    Span4Mux_v I__7522 (
            .O(N__38375),
            .I(N__38368));
    CEMux I__7521 (
            .O(N__38374),
            .I(N__38365));
    Odrv12 I__7520 (
            .O(N__38371),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__7519 (
            .O(N__38368),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    LocalMux I__7518 (
            .O(N__38365),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    CascadeMux I__7517 (
            .O(N__38358),
            .I(N__38355));
    InMux I__7516 (
            .O(N__38355),
            .I(N__38352));
    LocalMux I__7515 (
            .O(N__38352),
            .I(N__38349));
    Span4Mux_h I__7514 (
            .O(N__38349),
            .I(N__38346));
    Odrv4 I__7513 (
            .O(N__38346),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__7512 (
            .O(N__38343),
            .I(N__38338));
    InMux I__7511 (
            .O(N__38342),
            .I(N__38333));
    InMux I__7510 (
            .O(N__38341),
            .I(N__38333));
    LocalMux I__7509 (
            .O(N__38338),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ));
    LocalMux I__7508 (
            .O(N__38333),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ));
    InMux I__7507 (
            .O(N__38328),
            .I(N__38322));
    InMux I__7506 (
            .O(N__38327),
            .I(N__38322));
    LocalMux I__7505 (
            .O(N__38322),
            .I(N__38319));
    Span4Mux_v I__7504 (
            .O(N__38319),
            .I(N__38316));
    Odrv4 I__7503 (
            .O(N__38316),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ));
    CascadeMux I__7502 (
            .O(N__38313),
            .I(N__38309));
    InMux I__7501 (
            .O(N__38312),
            .I(N__38304));
    InMux I__7500 (
            .O(N__38309),
            .I(N__38304));
    LocalMux I__7499 (
            .O(N__38304),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ));
    CascadeMux I__7498 (
            .O(N__38301),
            .I(N__38296));
    InMux I__7497 (
            .O(N__38300),
            .I(N__38293));
    InMux I__7496 (
            .O(N__38299),
            .I(N__38288));
    InMux I__7495 (
            .O(N__38296),
            .I(N__38288));
    LocalMux I__7494 (
            .O(N__38293),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ));
    LocalMux I__7493 (
            .O(N__38288),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ));
    InMux I__7492 (
            .O(N__38283),
            .I(N__38280));
    LocalMux I__7491 (
            .O(N__38280),
            .I(N__38277));
    Span4Mux_h I__7490 (
            .O(N__38277),
            .I(N__38274));
    Odrv4 I__7489 (
            .O(N__38274),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt18 ));
    InMux I__7488 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__7487 (
            .O(N__38268),
            .I(N__38265));
    Span4Mux_s2_v I__7486 (
            .O(N__38265),
            .I(N__38262));
    Span4Mux_v I__7485 (
            .O(N__38262),
            .I(N__38257));
    InMux I__7484 (
            .O(N__38261),
            .I(N__38252));
    InMux I__7483 (
            .O(N__38260),
            .I(N__38252));
    Span4Mux_v I__7482 (
            .O(N__38257),
            .I(N__38247));
    LocalMux I__7481 (
            .O(N__38252),
            .I(N__38247));
    Span4Mux_v I__7480 (
            .O(N__38247),
            .I(N__38243));
    InMux I__7479 (
            .O(N__38246),
            .I(N__38240));
    Odrv4 I__7478 (
            .O(N__38243),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7477 (
            .O(N__38240),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__7476 (
            .O(N__38235),
            .I(N__38232));
    LocalMux I__7475 (
            .O(N__38232),
            .I(N__38229));
    Odrv12 I__7474 (
            .O(N__38229),
            .I(s2_phy_c));
    IoInMux I__7473 (
            .O(N__38226),
            .I(N__38223));
    LocalMux I__7472 (
            .O(N__38223),
            .I(\current_shift_inst.timer_s1.N_153_i ));
    CascadeMux I__7471 (
            .O(N__38220),
            .I(N__38216));
    InMux I__7470 (
            .O(N__38219),
            .I(N__38209));
    InMux I__7469 (
            .O(N__38216),
            .I(N__38206));
    InMux I__7468 (
            .O(N__38215),
            .I(N__38203));
    InMux I__7467 (
            .O(N__38214),
            .I(N__38200));
    InMux I__7466 (
            .O(N__38213),
            .I(N__38197));
    CascadeMux I__7465 (
            .O(N__38212),
            .I(N__38194));
    LocalMux I__7464 (
            .O(N__38209),
            .I(N__38191));
    LocalMux I__7463 (
            .O(N__38206),
            .I(N__38182));
    LocalMux I__7462 (
            .O(N__38203),
            .I(N__38182));
    LocalMux I__7461 (
            .O(N__38200),
            .I(N__38182));
    LocalMux I__7460 (
            .O(N__38197),
            .I(N__38182));
    InMux I__7459 (
            .O(N__38194),
            .I(N__38179));
    Span4Mux_h I__7458 (
            .O(N__38191),
            .I(N__38176));
    Odrv4 I__7457 (
            .O(N__38182),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__7456 (
            .O(N__38179),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7455 (
            .O(N__38176),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    CascadeMux I__7454 (
            .O(N__38169),
            .I(N__38166));
    InMux I__7453 (
            .O(N__38166),
            .I(N__38162));
    InMux I__7452 (
            .O(N__38165),
            .I(N__38159));
    LocalMux I__7451 (
            .O(N__38162),
            .I(N__38156));
    LocalMux I__7450 (
            .O(N__38159),
            .I(\phase_controller_inst2.stoper_hc.counter ));
    Odrv4 I__7449 (
            .O(N__38156),
            .I(\phase_controller_inst2.stoper_hc.counter ));
    InMux I__7448 (
            .O(N__38151),
            .I(N__38147));
    InMux I__7447 (
            .O(N__38150),
            .I(N__38144));
    LocalMux I__7446 (
            .O(N__38147),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ));
    LocalMux I__7445 (
            .O(N__38144),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ));
    InMux I__7444 (
            .O(N__38139),
            .I(N__38136));
    LocalMux I__7443 (
            .O(N__38136),
            .I(\phase_controller_inst2.stoper_hc.counter_i_0 ));
    InMux I__7442 (
            .O(N__38133),
            .I(N__38129));
    InMux I__7441 (
            .O(N__38132),
            .I(N__38126));
    LocalMux I__7440 (
            .O(N__38129),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ));
    LocalMux I__7439 (
            .O(N__38126),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ));
    InMux I__7438 (
            .O(N__38121),
            .I(N__38118));
    LocalMux I__7437 (
            .O(N__38118),
            .I(\phase_controller_inst2.stoper_hc.counter_i_1 ));
    InMux I__7436 (
            .O(N__38115),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__7435 (
            .O(N__38112),
            .I(bfn_13_26_0_));
    InMux I__7434 (
            .O(N__38109),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__7433 (
            .O(N__38106),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__7432 (
            .O(N__38103),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__7431 (
            .O(N__38100),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__7430 (
            .O(N__38097),
            .I(N__38067));
    InMux I__7429 (
            .O(N__38096),
            .I(N__38067));
    InMux I__7428 (
            .O(N__38095),
            .I(N__38058));
    InMux I__7427 (
            .O(N__38094),
            .I(N__38058));
    InMux I__7426 (
            .O(N__38093),
            .I(N__38058));
    InMux I__7425 (
            .O(N__38092),
            .I(N__38058));
    InMux I__7424 (
            .O(N__38091),
            .I(N__38045));
    InMux I__7423 (
            .O(N__38090),
            .I(N__38045));
    InMux I__7422 (
            .O(N__38089),
            .I(N__38045));
    InMux I__7421 (
            .O(N__38088),
            .I(N__38045));
    InMux I__7420 (
            .O(N__38087),
            .I(N__38036));
    InMux I__7419 (
            .O(N__38086),
            .I(N__38036));
    InMux I__7418 (
            .O(N__38085),
            .I(N__38036));
    InMux I__7417 (
            .O(N__38084),
            .I(N__38036));
    InMux I__7416 (
            .O(N__38083),
            .I(N__38027));
    InMux I__7415 (
            .O(N__38082),
            .I(N__38027));
    InMux I__7414 (
            .O(N__38081),
            .I(N__38027));
    InMux I__7413 (
            .O(N__38080),
            .I(N__38027));
    InMux I__7412 (
            .O(N__38079),
            .I(N__38018));
    InMux I__7411 (
            .O(N__38078),
            .I(N__38018));
    InMux I__7410 (
            .O(N__38077),
            .I(N__38018));
    InMux I__7409 (
            .O(N__38076),
            .I(N__38018));
    InMux I__7408 (
            .O(N__38075),
            .I(N__38009));
    InMux I__7407 (
            .O(N__38074),
            .I(N__38009));
    InMux I__7406 (
            .O(N__38073),
            .I(N__38009));
    InMux I__7405 (
            .O(N__38072),
            .I(N__38009));
    LocalMux I__7404 (
            .O(N__38067),
            .I(N__38004));
    LocalMux I__7403 (
            .O(N__38058),
            .I(N__38004));
    InMux I__7402 (
            .O(N__38057),
            .I(N__37995));
    InMux I__7401 (
            .O(N__38056),
            .I(N__37995));
    InMux I__7400 (
            .O(N__38055),
            .I(N__37995));
    InMux I__7399 (
            .O(N__38054),
            .I(N__37995));
    LocalMux I__7398 (
            .O(N__38045),
            .I(N__37982));
    LocalMux I__7397 (
            .O(N__38036),
            .I(N__37982));
    LocalMux I__7396 (
            .O(N__38027),
            .I(N__37982));
    LocalMux I__7395 (
            .O(N__38018),
            .I(N__37982));
    LocalMux I__7394 (
            .O(N__38009),
            .I(N__37982));
    Span4Mux_v I__7393 (
            .O(N__38004),
            .I(N__37982));
    LocalMux I__7392 (
            .O(N__37995),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__7391 (
            .O(N__37982),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__7390 (
            .O(N__37977),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__7389 (
            .O(N__37974),
            .I(N__37969));
    CEMux I__7388 (
            .O(N__37973),
            .I(N__37965));
    CEMux I__7387 (
            .O(N__37972),
            .I(N__37962));
    LocalMux I__7386 (
            .O(N__37969),
            .I(N__37959));
    CEMux I__7385 (
            .O(N__37968),
            .I(N__37956));
    LocalMux I__7384 (
            .O(N__37965),
            .I(N__37951));
    LocalMux I__7383 (
            .O(N__37962),
            .I(N__37951));
    Span4Mux_v I__7382 (
            .O(N__37959),
            .I(N__37946));
    LocalMux I__7381 (
            .O(N__37956),
            .I(N__37946));
    Span4Mux_v I__7380 (
            .O(N__37951),
            .I(N__37943));
    Span4Mux_v I__7379 (
            .O(N__37946),
            .I(N__37940));
    Span4Mux_h I__7378 (
            .O(N__37943),
            .I(N__37937));
    Odrv4 I__7377 (
            .O(N__37940),
            .I(\delay_measurement_inst.delay_tr_timer.N_158_i ));
    Odrv4 I__7376 (
            .O(N__37937),
            .I(\delay_measurement_inst.delay_tr_timer.N_158_i ));
    InMux I__7375 (
            .O(N__37932),
            .I(N__37929));
    LocalMux I__7374 (
            .O(N__37929),
            .I(N__37926));
    Odrv4 I__7373 (
            .O(N__37926),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt16 ));
    InMux I__7372 (
            .O(N__37923),
            .I(N__37916));
    InMux I__7371 (
            .O(N__37922),
            .I(N__37916));
    InMux I__7370 (
            .O(N__37921),
            .I(N__37913));
    LocalMux I__7369 (
            .O(N__37916),
            .I(N__37910));
    LocalMux I__7368 (
            .O(N__37913),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    Odrv4 I__7367 (
            .O(N__37910),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    InMux I__7366 (
            .O(N__37905),
            .I(N__37899));
    InMux I__7365 (
            .O(N__37904),
            .I(N__37899));
    LocalMux I__7364 (
            .O(N__37899),
            .I(N__37896));
    Span4Mux_v I__7363 (
            .O(N__37896),
            .I(N__37893));
    Odrv4 I__7362 (
            .O(N__37893),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ));
    CascadeMux I__7361 (
            .O(N__37890),
            .I(N__37886));
    CascadeMux I__7360 (
            .O(N__37889),
            .I(N__37883));
    InMux I__7359 (
            .O(N__37886),
            .I(N__37878));
    InMux I__7358 (
            .O(N__37883),
            .I(N__37878));
    LocalMux I__7357 (
            .O(N__37878),
            .I(N__37875));
    Span4Mux_v I__7356 (
            .O(N__37875),
            .I(N__37872));
    Odrv4 I__7355 (
            .O(N__37872),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ));
    InMux I__7354 (
            .O(N__37869),
            .I(N__37862));
    InMux I__7353 (
            .O(N__37868),
            .I(N__37862));
    InMux I__7352 (
            .O(N__37867),
            .I(N__37859));
    LocalMux I__7351 (
            .O(N__37862),
            .I(N__37856));
    LocalMux I__7350 (
            .O(N__37859),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    Odrv4 I__7349 (
            .O(N__37856),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    CascadeMux I__7348 (
            .O(N__37851),
            .I(N__37848));
    InMux I__7347 (
            .O(N__37848),
            .I(N__37845));
    LocalMux I__7346 (
            .O(N__37845),
            .I(N__37842));
    Odrv4 I__7345 (
            .O(N__37842),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__7344 (
            .O(N__37839),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__7343 (
            .O(N__37836),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__7342 (
            .O(N__37833),
            .I(bfn_13_25_0_));
    InMux I__7341 (
            .O(N__37830),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__7340 (
            .O(N__37827),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__7339 (
            .O(N__37824),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__7338 (
            .O(N__37821),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__7337 (
            .O(N__37818),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__7336 (
            .O(N__37815),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__7335 (
            .O(N__37812),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__7334 (
            .O(N__37809),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__7333 (
            .O(N__37806),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__7332 (
            .O(N__37803),
            .I(bfn_13_24_0_));
    InMux I__7331 (
            .O(N__37800),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__7330 (
            .O(N__37797),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__7329 (
            .O(N__37794),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__7328 (
            .O(N__37791),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__7327 (
            .O(N__37788),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__7326 (
            .O(N__37785),
            .I(N__37782));
    LocalMux I__7325 (
            .O(N__37782),
            .I(N__37779));
    Span12Mux_v I__7324 (
            .O(N__37779),
            .I(N__37775));
    InMux I__7323 (
            .O(N__37778),
            .I(N__37772));
    Odrv12 I__7322 (
            .O(N__37775),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_26));
    LocalMux I__7321 (
            .O(N__37772),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_26));
    InMux I__7320 (
            .O(N__37767),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ));
    InMux I__7319 (
            .O(N__37764),
            .I(N__37761));
    LocalMux I__7318 (
            .O(N__37761),
            .I(N__37758));
    Span12Mux_v I__7317 (
            .O(N__37758),
            .I(N__37754));
    InMux I__7316 (
            .O(N__37757),
            .I(N__37751));
    Odrv12 I__7315 (
            .O(N__37754),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_27));
    LocalMux I__7314 (
            .O(N__37751),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_27));
    InMux I__7313 (
            .O(N__37746),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ));
    InMux I__7312 (
            .O(N__37743),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ));
    InMux I__7311 (
            .O(N__37740),
            .I(N__37734));
    InMux I__7310 (
            .O(N__37739),
            .I(N__37731));
    InMux I__7309 (
            .O(N__37738),
            .I(N__37728));
    InMux I__7308 (
            .O(N__37737),
            .I(N__37725));
    LocalMux I__7307 (
            .O(N__37734),
            .I(N__37720));
    LocalMux I__7306 (
            .O(N__37731),
            .I(N__37720));
    LocalMux I__7305 (
            .O(N__37728),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__7304 (
            .O(N__37725),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__7303 (
            .O(N__37720),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__7302 (
            .O(N__37713),
            .I(bfn_13_23_0_));
    InMux I__7301 (
            .O(N__37710),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__7300 (
            .O(N__37707),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__7299 (
            .O(N__37704),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__7298 (
            .O(N__37701),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__7297 (
            .O(N__37698),
            .I(N__37695));
    LocalMux I__7296 (
            .O(N__37695),
            .I(N__37691));
    InMux I__7295 (
            .O(N__37694),
            .I(N__37688));
    Odrv12 I__7294 (
            .O(N__37691),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_18));
    LocalMux I__7293 (
            .O(N__37688),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_18));
    InMux I__7292 (
            .O(N__37683),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ));
    InMux I__7291 (
            .O(N__37680),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ));
    InMux I__7290 (
            .O(N__37677),
            .I(N__37673));
    InMux I__7289 (
            .O(N__37676),
            .I(N__37670));
    LocalMux I__7288 (
            .O(N__37673),
            .I(N__37667));
    LocalMux I__7287 (
            .O(N__37670),
            .I(N__37664));
    Sp12to4 I__7286 (
            .O(N__37667),
            .I(N__37661));
    Odrv4 I__7285 (
            .O(N__37664),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_20));
    Odrv12 I__7284 (
            .O(N__37661),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_20));
    InMux I__7283 (
            .O(N__37656),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ));
    InMux I__7282 (
            .O(N__37653),
            .I(N__37650));
    LocalMux I__7281 (
            .O(N__37650),
            .I(N__37647));
    Span12Mux_v I__7280 (
            .O(N__37647),
            .I(N__37643));
    InMux I__7279 (
            .O(N__37646),
            .I(N__37640));
    Odrv12 I__7278 (
            .O(N__37643),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_21));
    LocalMux I__7277 (
            .O(N__37640),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_21));
    InMux I__7276 (
            .O(N__37635),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ));
    InMux I__7275 (
            .O(N__37632),
            .I(N__37629));
    LocalMux I__7274 (
            .O(N__37629),
            .I(N__37626));
    Span12Mux_v I__7273 (
            .O(N__37626),
            .I(N__37622));
    InMux I__7272 (
            .O(N__37625),
            .I(N__37619));
    Odrv12 I__7271 (
            .O(N__37622),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_22));
    LocalMux I__7270 (
            .O(N__37619),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_22));
    InMux I__7269 (
            .O(N__37614),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ));
    InMux I__7268 (
            .O(N__37611),
            .I(N__37608));
    LocalMux I__7267 (
            .O(N__37608),
            .I(N__37605));
    Span12Mux_v I__7266 (
            .O(N__37605),
            .I(N__37601));
    InMux I__7265 (
            .O(N__37604),
            .I(N__37598));
    Odrv12 I__7264 (
            .O(N__37601),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_23));
    LocalMux I__7263 (
            .O(N__37598),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_23));
    InMux I__7262 (
            .O(N__37593),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ));
    InMux I__7261 (
            .O(N__37590),
            .I(N__37587));
    LocalMux I__7260 (
            .O(N__37587),
            .I(N__37584));
    Sp12to4 I__7259 (
            .O(N__37584),
            .I(N__37580));
    InMux I__7258 (
            .O(N__37583),
            .I(N__37577));
    Odrv12 I__7257 (
            .O(N__37580),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_24));
    LocalMux I__7256 (
            .O(N__37577),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_24));
    InMux I__7255 (
            .O(N__37572),
            .I(bfn_13_22_0_));
    InMux I__7254 (
            .O(N__37569),
            .I(N__37566));
    LocalMux I__7253 (
            .O(N__37566),
            .I(N__37563));
    Sp12to4 I__7252 (
            .O(N__37563),
            .I(N__37559));
    InMux I__7251 (
            .O(N__37562),
            .I(N__37556));
    Odrv12 I__7250 (
            .O(N__37559),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_25));
    LocalMux I__7249 (
            .O(N__37556),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_25));
    InMux I__7248 (
            .O(N__37551),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ));
    InMux I__7247 (
            .O(N__37548),
            .I(N__37545));
    LocalMux I__7246 (
            .O(N__37545),
            .I(N__37542));
    Span4Mux_v I__7245 (
            .O(N__37542),
            .I(N__37538));
    InMux I__7244 (
            .O(N__37541),
            .I(N__37535));
    Span4Mux_v I__7243 (
            .O(N__37538),
            .I(N__37530));
    LocalMux I__7242 (
            .O(N__37535),
            .I(N__37530));
    Odrv4 I__7241 (
            .O(N__37530),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_9));
    InMux I__7240 (
            .O(N__37527),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ));
    InMux I__7239 (
            .O(N__37524),
            .I(N__37521));
    LocalMux I__7238 (
            .O(N__37521),
            .I(N__37518));
    Span4Mux_v I__7237 (
            .O(N__37518),
            .I(N__37514));
    InMux I__7236 (
            .O(N__37517),
            .I(N__37511));
    Odrv4 I__7235 (
            .O(N__37514),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_10));
    LocalMux I__7234 (
            .O(N__37511),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_10));
    InMux I__7233 (
            .O(N__37506),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ));
    InMux I__7232 (
            .O(N__37503),
            .I(N__37500));
    LocalMux I__7231 (
            .O(N__37500),
            .I(N__37497));
    Span4Mux_v I__7230 (
            .O(N__37497),
            .I(N__37493));
    InMux I__7229 (
            .O(N__37496),
            .I(N__37490));
    Odrv4 I__7228 (
            .O(N__37493),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_11));
    LocalMux I__7227 (
            .O(N__37490),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_11));
    InMux I__7226 (
            .O(N__37485),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ));
    InMux I__7225 (
            .O(N__37482),
            .I(N__37479));
    LocalMux I__7224 (
            .O(N__37479),
            .I(N__37476));
    Span4Mux_v I__7223 (
            .O(N__37476),
            .I(N__37472));
    InMux I__7222 (
            .O(N__37475),
            .I(N__37469));
    Odrv4 I__7221 (
            .O(N__37472),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_12));
    LocalMux I__7220 (
            .O(N__37469),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_12));
    InMux I__7219 (
            .O(N__37464),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ));
    InMux I__7218 (
            .O(N__37461),
            .I(N__37458));
    LocalMux I__7217 (
            .O(N__37458),
            .I(N__37455));
    Span12Mux_v I__7216 (
            .O(N__37455),
            .I(N__37451));
    InMux I__7215 (
            .O(N__37454),
            .I(N__37448));
    Odrv12 I__7214 (
            .O(N__37451),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_13));
    LocalMux I__7213 (
            .O(N__37448),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_13));
    InMux I__7212 (
            .O(N__37443),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ));
    InMux I__7211 (
            .O(N__37440),
            .I(N__37437));
    LocalMux I__7210 (
            .O(N__37437),
            .I(N__37434));
    Span4Mux_v I__7209 (
            .O(N__37434),
            .I(N__37430));
    InMux I__7208 (
            .O(N__37433),
            .I(N__37427));
    Odrv4 I__7207 (
            .O(N__37430),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_14));
    LocalMux I__7206 (
            .O(N__37427),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_14));
    InMux I__7205 (
            .O(N__37422),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ));
    InMux I__7204 (
            .O(N__37419),
            .I(N__37416));
    LocalMux I__7203 (
            .O(N__37416),
            .I(N__37413));
    Span12Mux_v I__7202 (
            .O(N__37413),
            .I(N__37409));
    InMux I__7201 (
            .O(N__37412),
            .I(N__37406));
    Odrv12 I__7200 (
            .O(N__37409),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_15));
    LocalMux I__7199 (
            .O(N__37406),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_15));
    InMux I__7198 (
            .O(N__37401),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ));
    InMux I__7197 (
            .O(N__37398),
            .I(N__37395));
    LocalMux I__7196 (
            .O(N__37395),
            .I(N__37392));
    Span12Mux_v I__7195 (
            .O(N__37392),
            .I(N__37388));
    InMux I__7194 (
            .O(N__37391),
            .I(N__37385));
    Odrv12 I__7193 (
            .O(N__37388),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_16));
    LocalMux I__7192 (
            .O(N__37385),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_16));
    InMux I__7191 (
            .O(N__37380),
            .I(bfn_13_21_0_));
    InMux I__7190 (
            .O(N__37377),
            .I(N__37374));
    LocalMux I__7189 (
            .O(N__37374),
            .I(N__37370));
    InMux I__7188 (
            .O(N__37373),
            .I(N__37367));
    Sp12to4 I__7187 (
            .O(N__37370),
            .I(N__37364));
    LocalMux I__7186 (
            .O(N__37367),
            .I(N__37361));
    Odrv12 I__7185 (
            .O(N__37364),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_17));
    Odrv4 I__7184 (
            .O(N__37361),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_17));
    InMux I__7183 (
            .O(N__37356),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ));
    InMux I__7182 (
            .O(N__37353),
            .I(N__37349));
    InMux I__7181 (
            .O(N__37352),
            .I(N__37346));
    LocalMux I__7180 (
            .O(N__37349),
            .I(N__37343));
    LocalMux I__7179 (
            .O(N__37346),
            .I(N__37340));
    Sp12to4 I__7178 (
            .O(N__37343),
            .I(N__37337));
    Span4Mux_v I__7177 (
            .O(N__37340),
            .I(N__37334));
    Span12Mux_s7_v I__7176 (
            .O(N__37337),
            .I(N__37331));
    Odrv4 I__7175 (
            .O(N__37334),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_1));
    Odrv12 I__7174 (
            .O(N__37331),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_1));
    InMux I__7173 (
            .O(N__37326),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ));
    InMux I__7172 (
            .O(N__37323),
            .I(N__37320));
    LocalMux I__7171 (
            .O(N__37320),
            .I(N__37316));
    InMux I__7170 (
            .O(N__37319),
            .I(N__37313));
    Span12Mux_h I__7169 (
            .O(N__37316),
            .I(N__37310));
    LocalMux I__7168 (
            .O(N__37313),
            .I(N__37307));
    Span12Mux_v I__7167 (
            .O(N__37310),
            .I(N__37304));
    Span4Mux_v I__7166 (
            .O(N__37307),
            .I(N__37301));
    Odrv12 I__7165 (
            .O(N__37304),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_2));
    Odrv4 I__7164 (
            .O(N__37301),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_2));
    InMux I__7163 (
            .O(N__37296),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ));
    InMux I__7162 (
            .O(N__37293),
            .I(N__37290));
    LocalMux I__7161 (
            .O(N__37290),
            .I(N__37286));
    InMux I__7160 (
            .O(N__37289),
            .I(N__37283));
    Sp12to4 I__7159 (
            .O(N__37286),
            .I(N__37280));
    LocalMux I__7158 (
            .O(N__37283),
            .I(N__37277));
    Span12Mux_v I__7157 (
            .O(N__37280),
            .I(N__37274));
    Span4Mux_v I__7156 (
            .O(N__37277),
            .I(N__37271));
    Odrv12 I__7155 (
            .O(N__37274),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_3));
    Odrv4 I__7154 (
            .O(N__37271),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_3));
    InMux I__7153 (
            .O(N__37266),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ));
    InMux I__7152 (
            .O(N__37263),
            .I(N__37259));
    InMux I__7151 (
            .O(N__37262),
            .I(N__37256));
    LocalMux I__7150 (
            .O(N__37259),
            .I(N__37253));
    LocalMux I__7149 (
            .O(N__37256),
            .I(N__37250));
    Span4Mux_h I__7148 (
            .O(N__37253),
            .I(N__37247));
    Span4Mux_v I__7147 (
            .O(N__37250),
            .I(N__37244));
    Span4Mux_v I__7146 (
            .O(N__37247),
            .I(N__37241));
    Odrv4 I__7145 (
            .O(N__37244),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_4));
    Odrv4 I__7144 (
            .O(N__37241),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_4));
    InMux I__7143 (
            .O(N__37236),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ));
    InMux I__7142 (
            .O(N__37233),
            .I(N__37230));
    LocalMux I__7141 (
            .O(N__37230),
            .I(N__37226));
    InMux I__7140 (
            .O(N__37229),
            .I(N__37223));
    Span12Mux_s6_v I__7139 (
            .O(N__37226),
            .I(N__37220));
    LocalMux I__7138 (
            .O(N__37223),
            .I(N__37217));
    Span12Mux_v I__7137 (
            .O(N__37220),
            .I(N__37214));
    Span4Mux_v I__7136 (
            .O(N__37217),
            .I(N__37211));
    Odrv12 I__7135 (
            .O(N__37214),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_5));
    Odrv4 I__7134 (
            .O(N__37211),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_5));
    InMux I__7133 (
            .O(N__37206),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ));
    InMux I__7132 (
            .O(N__37203),
            .I(N__37199));
    InMux I__7131 (
            .O(N__37202),
            .I(N__37196));
    LocalMux I__7130 (
            .O(N__37199),
            .I(N__37193));
    LocalMux I__7129 (
            .O(N__37196),
            .I(N__37190));
    Span4Mux_v I__7128 (
            .O(N__37193),
            .I(N__37187));
    Span4Mux_v I__7127 (
            .O(N__37190),
            .I(N__37184));
    Odrv4 I__7126 (
            .O(N__37187),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_6));
    Odrv4 I__7125 (
            .O(N__37184),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_6));
    InMux I__7124 (
            .O(N__37179),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ));
    InMux I__7123 (
            .O(N__37176),
            .I(N__37173));
    LocalMux I__7122 (
            .O(N__37173),
            .I(N__37169));
    InMux I__7121 (
            .O(N__37172),
            .I(N__37166));
    Span4Mux_v I__7120 (
            .O(N__37169),
            .I(N__37163));
    LocalMux I__7119 (
            .O(N__37166),
            .I(N__37160));
    Odrv4 I__7118 (
            .O(N__37163),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_7));
    Odrv4 I__7117 (
            .O(N__37160),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_7));
    InMux I__7116 (
            .O(N__37155),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ));
    InMux I__7115 (
            .O(N__37152),
            .I(N__37149));
    LocalMux I__7114 (
            .O(N__37149),
            .I(N__37145));
    InMux I__7113 (
            .O(N__37148),
            .I(N__37142));
    Sp12to4 I__7112 (
            .O(N__37145),
            .I(N__37139));
    LocalMux I__7111 (
            .O(N__37142),
            .I(N__37136));
    Span12Mux_v I__7110 (
            .O(N__37139),
            .I(N__37133));
    Span4Mux_v I__7109 (
            .O(N__37136),
            .I(N__37130));
    Odrv12 I__7108 (
            .O(N__37133),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_8));
    Odrv4 I__7107 (
            .O(N__37130),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_8));
    InMux I__7106 (
            .O(N__37125),
            .I(bfn_13_20_0_));
    InMux I__7105 (
            .O(N__37122),
            .I(N__37119));
    LocalMux I__7104 (
            .O(N__37119),
            .I(N__37116));
    Span4Mux_v I__7103 (
            .O(N__37116),
            .I(N__37113));
    Span4Mux_h I__7102 (
            .O(N__37113),
            .I(N__37110));
    Odrv4 I__7101 (
            .O(N__37110),
            .I(\phase_controller_inst1.stoper_tr.un4_start_0 ));
    CascadeMux I__7100 (
            .O(N__37107),
            .I(N__37103));
    InMux I__7099 (
            .O(N__37106),
            .I(N__37095));
    InMux I__7098 (
            .O(N__37103),
            .I(N__37095));
    InMux I__7097 (
            .O(N__37102),
            .I(N__37095));
    LocalMux I__7096 (
            .O(N__37095),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__7095 (
            .O(N__37092),
            .I(N__37086));
    InMux I__7094 (
            .O(N__37091),
            .I(N__37086));
    LocalMux I__7093 (
            .O(N__37086),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CascadeMux I__7092 (
            .O(N__37083),
            .I(N__37079));
    InMux I__7091 (
            .O(N__37082),
            .I(N__37076));
    InMux I__7090 (
            .O(N__37079),
            .I(N__37073));
    LocalMux I__7089 (
            .O(N__37076),
            .I(N__37067));
    LocalMux I__7088 (
            .O(N__37073),
            .I(N__37067));
    InMux I__7087 (
            .O(N__37072),
            .I(N__37064));
    Span4Mux_v I__7086 (
            .O(N__37067),
            .I(N__37059));
    LocalMux I__7085 (
            .O(N__37064),
            .I(N__37059));
    Span4Mux_h I__7084 (
            .O(N__37059),
            .I(N__37056));
    Sp12to4 I__7083 (
            .O(N__37056),
            .I(N__37053));
    Span12Mux_v I__7082 (
            .O(N__37053),
            .I(N__37050));
    Odrv12 I__7081 (
            .O(N__37050),
            .I(il_min_comp1_c));
    InMux I__7080 (
            .O(N__37047),
            .I(N__37044));
    LocalMux I__7079 (
            .O(N__37044),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__7078 (
            .O(N__37041),
            .I(N__37037));
    InMux I__7077 (
            .O(N__37040),
            .I(N__37033));
    LocalMux I__7076 (
            .O(N__37037),
            .I(N__37028));
    InMux I__7075 (
            .O(N__37036),
            .I(N__37025));
    LocalMux I__7074 (
            .O(N__37033),
            .I(N__37022));
    InMux I__7073 (
            .O(N__37032),
            .I(N__37017));
    InMux I__7072 (
            .O(N__37031),
            .I(N__37017));
    Span4Mux_v I__7071 (
            .O(N__37028),
            .I(N__37014));
    LocalMux I__7070 (
            .O(N__37025),
            .I(N__37010));
    Span4Mux_h I__7069 (
            .O(N__37022),
            .I(N__37007));
    LocalMux I__7068 (
            .O(N__37017),
            .I(N__37002));
    Span4Mux_h I__7067 (
            .O(N__37014),
            .I(N__37002));
    InMux I__7066 (
            .O(N__37013),
            .I(N__36999));
    Span4Mux_h I__7065 (
            .O(N__37010),
            .I(N__36996));
    Span4Mux_v I__7064 (
            .O(N__37007),
            .I(N__36993));
    Sp12to4 I__7063 (
            .O(N__37002),
            .I(N__36990));
    LocalMux I__7062 (
            .O(N__36999),
            .I(N__36985));
    Span4Mux_v I__7061 (
            .O(N__36996),
            .I(N__36985));
    Odrv4 I__7060 (
            .O(N__36993),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__7059 (
            .O(N__36990),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__7058 (
            .O(N__36985),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__7057 (
            .O(N__36978),
            .I(N__36975));
    InMux I__7056 (
            .O(N__36975),
            .I(N__36971));
    InMux I__7055 (
            .O(N__36974),
            .I(N__36967));
    LocalMux I__7054 (
            .O(N__36971),
            .I(N__36963));
    InMux I__7053 (
            .O(N__36970),
            .I(N__36960));
    LocalMux I__7052 (
            .O(N__36967),
            .I(N__36956));
    InMux I__7051 (
            .O(N__36966),
            .I(N__36953));
    Span4Mux_h I__7050 (
            .O(N__36963),
            .I(N__36950));
    LocalMux I__7049 (
            .O(N__36960),
            .I(N__36946));
    InMux I__7048 (
            .O(N__36959),
            .I(N__36943));
    Span4Mux_h I__7047 (
            .O(N__36956),
            .I(N__36940));
    LocalMux I__7046 (
            .O(N__36953),
            .I(N__36937));
    Span4Mux_v I__7045 (
            .O(N__36950),
            .I(N__36934));
    InMux I__7044 (
            .O(N__36949),
            .I(N__36931));
    Span12Mux_v I__7043 (
            .O(N__36946),
            .I(N__36928));
    LocalMux I__7042 (
            .O(N__36943),
            .I(N__36921));
    Span4Mux_v I__7041 (
            .O(N__36940),
            .I(N__36921));
    Span4Mux_s3_v I__7040 (
            .O(N__36937),
            .I(N__36921));
    Odrv4 I__7039 (
            .O(N__36934),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__7038 (
            .O(N__36931),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv12 I__7037 (
            .O(N__36928),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__7036 (
            .O(N__36921),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__7035 (
            .O(N__36912),
            .I(N__36906));
    InMux I__7034 (
            .O(N__36911),
            .I(N__36906));
    LocalMux I__7033 (
            .O(N__36906),
            .I(N__36903));
    Span4Mux_h I__7032 (
            .O(N__36903),
            .I(N__36900));
    Span4Mux_v I__7031 (
            .O(N__36900),
            .I(N__36897));
    Span4Mux_v I__7030 (
            .O(N__36897),
            .I(N__36893));
    InMux I__7029 (
            .O(N__36896),
            .I(N__36890));
    Odrv4 I__7028 (
            .O(N__36893),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ));
    LocalMux I__7027 (
            .O(N__36890),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ));
    InMux I__7026 (
            .O(N__36885),
            .I(N__36882));
    LocalMux I__7025 (
            .O(N__36882),
            .I(N__36878));
    CascadeMux I__7024 (
            .O(N__36881),
            .I(N__36874));
    Span4Mux_h I__7023 (
            .O(N__36878),
            .I(N__36871));
    InMux I__7022 (
            .O(N__36877),
            .I(N__36866));
    InMux I__7021 (
            .O(N__36874),
            .I(N__36866));
    Span4Mux_v I__7020 (
            .O(N__36871),
            .I(N__36863));
    LocalMux I__7019 (
            .O(N__36866),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    Odrv4 I__7018 (
            .O(N__36863),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    CascadeMux I__7017 (
            .O(N__36858),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__7016 (
            .O(N__36855),
            .I(N__36852));
    LocalMux I__7015 (
            .O(N__36852),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    CascadeMux I__7014 (
            .O(N__36849),
            .I(N__36846));
    InMux I__7013 (
            .O(N__36846),
            .I(N__36840));
    InMux I__7012 (
            .O(N__36845),
            .I(N__36835));
    InMux I__7011 (
            .O(N__36844),
            .I(N__36835));
    InMux I__7010 (
            .O(N__36843),
            .I(N__36832));
    LocalMux I__7009 (
            .O(N__36840),
            .I(N__36829));
    LocalMux I__7008 (
            .O(N__36835),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__7007 (
            .O(N__36832),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__7006 (
            .O(N__36829),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__7005 (
            .O(N__36822),
            .I(N__36818));
    InMux I__7004 (
            .O(N__36821),
            .I(N__36814));
    LocalMux I__7003 (
            .O(N__36818),
            .I(N__36811));
    InMux I__7002 (
            .O(N__36817),
            .I(N__36808));
    LocalMux I__7001 (
            .O(N__36814),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__7000 (
            .O(N__36811),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__6999 (
            .O(N__36808),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__6998 (
            .O(N__36801),
            .I(N__36798));
    LocalMux I__6997 (
            .O(N__36798),
            .I(\phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ));
    InMux I__6996 (
            .O(N__36795),
            .I(N__36791));
    InMux I__6995 (
            .O(N__36794),
            .I(N__36788));
    LocalMux I__6994 (
            .O(N__36791),
            .I(N__36784));
    LocalMux I__6993 (
            .O(N__36788),
            .I(N__36780));
    InMux I__6992 (
            .O(N__36787),
            .I(N__36777));
    Span4Mux_h I__6991 (
            .O(N__36784),
            .I(N__36774));
    InMux I__6990 (
            .O(N__36783),
            .I(N__36771));
    Span4Mux_v I__6989 (
            .O(N__36780),
            .I(N__36768));
    LocalMux I__6988 (
            .O(N__36777),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__6987 (
            .O(N__36774),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__6986 (
            .O(N__36771),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__6985 (
            .O(N__36768),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__6984 (
            .O(N__36759),
            .I(N__36755));
    CascadeMux I__6983 (
            .O(N__36758),
            .I(N__36750));
    LocalMux I__6982 (
            .O(N__36755),
            .I(N__36747));
    InMux I__6981 (
            .O(N__36754),
            .I(N__36744));
    InMux I__6980 (
            .O(N__36753),
            .I(N__36739));
    InMux I__6979 (
            .O(N__36750),
            .I(N__36739));
    Span4Mux_v I__6978 (
            .O(N__36747),
            .I(N__36736));
    LocalMux I__6977 (
            .O(N__36744),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6976 (
            .O(N__36739),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__6975 (
            .O(N__36736),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__6974 (
            .O(N__36729),
            .I(N__36725));
    InMux I__6973 (
            .O(N__36728),
            .I(N__36722));
    LocalMux I__6972 (
            .O(N__36725),
            .I(N__36719));
    LocalMux I__6971 (
            .O(N__36722),
            .I(N__36716));
    Span12Mux_v I__6970 (
            .O(N__36719),
            .I(N__36713));
    Odrv12 I__6969 (
            .O(N__36716),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv12 I__6968 (
            .O(N__36713),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__6967 (
            .O(N__36708),
            .I(N__36704));
    InMux I__6966 (
            .O(N__36707),
            .I(N__36701));
    InMux I__6965 (
            .O(N__36704),
            .I(N__36698));
    LocalMux I__6964 (
            .O(N__36701),
            .I(N__36694));
    LocalMux I__6963 (
            .O(N__36698),
            .I(N__36691));
    CascadeMux I__6962 (
            .O(N__36697),
            .I(N__36688));
    Span4Mux_v I__6961 (
            .O(N__36694),
            .I(N__36685));
    Span4Mux_v I__6960 (
            .O(N__36691),
            .I(N__36682));
    InMux I__6959 (
            .O(N__36688),
            .I(N__36678));
    Sp12to4 I__6958 (
            .O(N__36685),
            .I(N__36673));
    Sp12to4 I__6957 (
            .O(N__36682),
            .I(N__36673));
    InMux I__6956 (
            .O(N__36681),
            .I(N__36670));
    LocalMux I__6955 (
            .O(N__36678),
            .I(N__36667));
    Span12Mux_h I__6954 (
            .O(N__36673),
            .I(N__36664));
    LocalMux I__6953 (
            .O(N__36670),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__6952 (
            .O(N__36667),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__6951 (
            .O(N__36664),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__6950 (
            .O(N__36657),
            .I(N__36654));
    LocalMux I__6949 (
            .O(N__36654),
            .I(N__36650));
    InMux I__6948 (
            .O(N__36653),
            .I(N__36647));
    Span4Mux_h I__6947 (
            .O(N__36650),
            .I(N__36641));
    LocalMux I__6946 (
            .O(N__36647),
            .I(N__36641));
    InMux I__6945 (
            .O(N__36646),
            .I(N__36638));
    Span4Mux_v I__6944 (
            .O(N__36641),
            .I(N__36635));
    LocalMux I__6943 (
            .O(N__36638),
            .I(N__36632));
    Span4Mux_v I__6942 (
            .O(N__36635),
            .I(N__36629));
    Span4Mux_v I__6941 (
            .O(N__36632),
            .I(N__36626));
    Sp12to4 I__6940 (
            .O(N__36629),
            .I(N__36623));
    Span4Mux_h I__6939 (
            .O(N__36626),
            .I(N__36620));
    Span12Mux_h I__6938 (
            .O(N__36623),
            .I(N__36615));
    Sp12to4 I__6937 (
            .O(N__36620),
            .I(N__36615));
    Odrv12 I__6936 (
            .O(N__36615),
            .I(il_max_comp1_c));
    InMux I__6935 (
            .O(N__36612),
            .I(N__36608));
    InMux I__6934 (
            .O(N__36611),
            .I(N__36605));
    LocalMux I__6933 (
            .O(N__36608),
            .I(N__36601));
    LocalMux I__6932 (
            .O(N__36605),
            .I(N__36598));
    InMux I__6931 (
            .O(N__36604),
            .I(N__36595));
    Span4Mux_s3_v I__6930 (
            .O(N__36601),
            .I(N__36590));
    Span4Mux_s3_v I__6929 (
            .O(N__36598),
            .I(N__36590));
    LocalMux I__6928 (
            .O(N__36595),
            .I(N__36585));
    Span4Mux_h I__6927 (
            .O(N__36590),
            .I(N__36582));
    InMux I__6926 (
            .O(N__36589),
            .I(N__36577));
    InMux I__6925 (
            .O(N__36588),
            .I(N__36577));
    Span4Mux_v I__6924 (
            .O(N__36585),
            .I(N__36574));
    Sp12to4 I__6923 (
            .O(N__36582),
            .I(N__36571));
    LocalMux I__6922 (
            .O(N__36577),
            .I(N__36568));
    Span4Mux_h I__6921 (
            .O(N__36574),
            .I(N__36562));
    Span12Mux_s11_v I__6920 (
            .O(N__36571),
            .I(N__36557));
    Sp12to4 I__6919 (
            .O(N__36568),
            .I(N__36557));
    InMux I__6918 (
            .O(N__36567),
            .I(N__36550));
    InMux I__6917 (
            .O(N__36566),
            .I(N__36550));
    InMux I__6916 (
            .O(N__36565),
            .I(N__36550));
    Sp12to4 I__6915 (
            .O(N__36562),
            .I(N__36547));
    Span12Mux_v I__6914 (
            .O(N__36557),
            .I(N__36542));
    LocalMux I__6913 (
            .O(N__36550),
            .I(N__36542));
    Span12Mux_v I__6912 (
            .O(N__36547),
            .I(N__36537));
    Span12Mux_h I__6911 (
            .O(N__36542),
            .I(N__36537));
    Odrv12 I__6910 (
            .O(N__36537),
            .I(start_stop_c));
    InMux I__6909 (
            .O(N__36534),
            .I(N__36531));
    LocalMux I__6908 (
            .O(N__36531),
            .I(N__36526));
    InMux I__6907 (
            .O(N__36530),
            .I(N__36521));
    InMux I__6906 (
            .O(N__36529),
            .I(N__36521));
    Odrv12 I__6905 (
            .O(N__36526),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__6904 (
            .O(N__36521),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    CascadeMux I__6903 (
            .O(N__36516),
            .I(\phase_controller_inst1.state_ns_0_0_1_cascade_ ));
    InMux I__6902 (
            .O(N__36513),
            .I(N__36509));
    CascadeMux I__6901 (
            .O(N__36512),
            .I(N__36506));
    LocalMux I__6900 (
            .O(N__36509),
            .I(N__36502));
    InMux I__6899 (
            .O(N__36506),
            .I(N__36497));
    InMux I__6898 (
            .O(N__36505),
            .I(N__36497));
    Span12Mux_h I__6897 (
            .O(N__36502),
            .I(N__36494));
    LocalMux I__6896 (
            .O(N__36497),
            .I(\phase_controller_inst1.start_flagZ0 ));
    Odrv12 I__6895 (
            .O(N__36494),
            .I(\phase_controller_inst1.start_flagZ0 ));
    InMux I__6894 (
            .O(N__36489),
            .I(N__36486));
    LocalMux I__6893 (
            .O(N__36486),
            .I(N__36483));
    Span4Mux_h I__6892 (
            .O(N__36483),
            .I(N__36480));
    Odrv4 I__6891 (
            .O(N__36480),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ));
    InMux I__6890 (
            .O(N__36477),
            .I(N__36473));
    InMux I__6889 (
            .O(N__36476),
            .I(N__36470));
    LocalMux I__6888 (
            .O(N__36473),
            .I(N__36467));
    LocalMux I__6887 (
            .O(N__36470),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ));
    Odrv4 I__6886 (
            .O(N__36467),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ));
    InMux I__6885 (
            .O(N__36462),
            .I(N__36456));
    InMux I__6884 (
            .O(N__36461),
            .I(N__36456));
    LocalMux I__6883 (
            .O(N__36456),
            .I(N__36453));
    Span4Mux_h I__6882 (
            .O(N__36453),
            .I(N__36450));
    Odrv4 I__6881 (
            .O(N__36450),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ));
    CascadeMux I__6880 (
            .O(N__36447),
            .I(N__36443));
    CascadeMux I__6879 (
            .O(N__36446),
            .I(N__36440));
    InMux I__6878 (
            .O(N__36443),
            .I(N__36435));
    InMux I__6877 (
            .O(N__36440),
            .I(N__36435));
    LocalMux I__6876 (
            .O(N__36435),
            .I(N__36432));
    Span4Mux_h I__6875 (
            .O(N__36432),
            .I(N__36429));
    Odrv4 I__6874 (
            .O(N__36429),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ));
    InMux I__6873 (
            .O(N__36426),
            .I(N__36423));
    LocalMux I__6872 (
            .O(N__36423),
            .I(N__36420));
    Span4Mux_v I__6871 (
            .O(N__36420),
            .I(N__36417));
    Span4Mux_v I__6870 (
            .O(N__36417),
            .I(N__36414));
    Odrv4 I__6869 (
            .O(N__36414),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ));
    CascadeMux I__6868 (
            .O(N__36411),
            .I(N__36408));
    InMux I__6867 (
            .O(N__36408),
            .I(N__36402));
    InMux I__6866 (
            .O(N__36407),
            .I(N__36402));
    LocalMux I__6865 (
            .O(N__36402),
            .I(N__36399));
    Span4Mux_h I__6864 (
            .O(N__36399),
            .I(N__36396));
    Odrv4 I__6863 (
            .O(N__36396),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ));
    InMux I__6862 (
            .O(N__36393),
            .I(N__36387));
    InMux I__6861 (
            .O(N__36392),
            .I(N__36387));
    LocalMux I__6860 (
            .O(N__36387),
            .I(N__36384));
    Span4Mux_h I__6859 (
            .O(N__36384),
            .I(N__36381));
    Odrv4 I__6858 (
            .O(N__36381),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ));
    CascadeMux I__6857 (
            .O(N__36378),
            .I(N__36374));
    InMux I__6856 (
            .O(N__36377),
            .I(N__36369));
    InMux I__6855 (
            .O(N__36374),
            .I(N__36369));
    LocalMux I__6854 (
            .O(N__36369),
            .I(N__36366));
    Span4Mux_h I__6853 (
            .O(N__36366),
            .I(N__36363));
    Odrv4 I__6852 (
            .O(N__36363),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ));
    CascadeMux I__6851 (
            .O(N__36360),
            .I(N__36356));
    CascadeMux I__6850 (
            .O(N__36359),
            .I(N__36353));
    InMux I__6849 (
            .O(N__36356),
            .I(N__36348));
    InMux I__6848 (
            .O(N__36353),
            .I(N__36348));
    LocalMux I__6847 (
            .O(N__36348),
            .I(N__36345));
    Span4Mux_v I__6846 (
            .O(N__36345),
            .I(N__36342));
    Odrv4 I__6845 (
            .O(N__36342),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ));
    CEMux I__6844 (
            .O(N__36339),
            .I(N__36336));
    LocalMux I__6843 (
            .O(N__36336),
            .I(N__36329));
    CEMux I__6842 (
            .O(N__36335),
            .I(N__36326));
    CEMux I__6841 (
            .O(N__36334),
            .I(N__36321));
    CEMux I__6840 (
            .O(N__36333),
            .I(N__36318));
    CEMux I__6839 (
            .O(N__36332),
            .I(N__36315));
    Span4Mux_h I__6838 (
            .O(N__36329),
            .I(N__36309));
    LocalMux I__6837 (
            .O(N__36326),
            .I(N__36309));
    CEMux I__6836 (
            .O(N__36325),
            .I(N__36306));
    CEMux I__6835 (
            .O(N__36324),
            .I(N__36303));
    LocalMux I__6834 (
            .O(N__36321),
            .I(N__36298));
    LocalMux I__6833 (
            .O(N__36318),
            .I(N__36298));
    LocalMux I__6832 (
            .O(N__36315),
            .I(N__36295));
    CEMux I__6831 (
            .O(N__36314),
            .I(N__36292));
    Span4Mux_v I__6830 (
            .O(N__36309),
            .I(N__36289));
    LocalMux I__6829 (
            .O(N__36306),
            .I(N__36286));
    LocalMux I__6828 (
            .O(N__36303),
            .I(N__36283));
    Span4Mux_v I__6827 (
            .O(N__36298),
            .I(N__36276));
    Span4Mux_v I__6826 (
            .O(N__36295),
            .I(N__36276));
    LocalMux I__6825 (
            .O(N__36292),
            .I(N__36276));
    Span4Mux_h I__6824 (
            .O(N__36289),
            .I(N__36271));
    Span4Mux_v I__6823 (
            .O(N__36286),
            .I(N__36271));
    Span4Mux_v I__6822 (
            .O(N__36283),
            .I(N__36266));
    Span4Mux_v I__6821 (
            .O(N__36276),
            .I(N__36266));
    Odrv4 I__6820 (
            .O(N__36271),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__6819 (
            .O(N__36266),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    InMux I__6818 (
            .O(N__36261),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_25 ));
    InMux I__6817 (
            .O(N__36258),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_26 ));
    InMux I__6816 (
            .O(N__36255),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_27 ));
    InMux I__6815 (
            .O(N__36252),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_28 ));
    InMux I__6814 (
            .O(N__36249),
            .I(N__36244));
    InMux I__6813 (
            .O(N__36248),
            .I(N__36239));
    InMux I__6812 (
            .O(N__36247),
            .I(N__36239));
    LocalMux I__6811 (
            .O(N__36244),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    LocalMux I__6810 (
            .O(N__36239),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    InMux I__6809 (
            .O(N__36234),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_29 ));
    InMux I__6808 (
            .O(N__36231),
            .I(N__36214));
    InMux I__6807 (
            .O(N__36230),
            .I(N__36214));
    InMux I__6806 (
            .O(N__36229),
            .I(N__36214));
    InMux I__6805 (
            .O(N__36228),
            .I(N__36184));
    InMux I__6804 (
            .O(N__36227),
            .I(N__36184));
    InMux I__6803 (
            .O(N__36226),
            .I(N__36184));
    InMux I__6802 (
            .O(N__36225),
            .I(N__36184));
    InMux I__6801 (
            .O(N__36224),
            .I(N__36175));
    InMux I__6800 (
            .O(N__36223),
            .I(N__36175));
    InMux I__6799 (
            .O(N__36222),
            .I(N__36175));
    InMux I__6798 (
            .O(N__36221),
            .I(N__36175));
    LocalMux I__6797 (
            .O(N__36214),
            .I(N__36172));
    InMux I__6796 (
            .O(N__36213),
            .I(N__36163));
    InMux I__6795 (
            .O(N__36212),
            .I(N__36163));
    InMux I__6794 (
            .O(N__36211),
            .I(N__36163));
    InMux I__6793 (
            .O(N__36210),
            .I(N__36163));
    InMux I__6792 (
            .O(N__36209),
            .I(N__36154));
    InMux I__6791 (
            .O(N__36208),
            .I(N__36154));
    InMux I__6790 (
            .O(N__36207),
            .I(N__36154));
    InMux I__6789 (
            .O(N__36206),
            .I(N__36154));
    InMux I__6788 (
            .O(N__36205),
            .I(N__36145));
    InMux I__6787 (
            .O(N__36204),
            .I(N__36145));
    InMux I__6786 (
            .O(N__36203),
            .I(N__36145));
    InMux I__6785 (
            .O(N__36202),
            .I(N__36145));
    InMux I__6784 (
            .O(N__36201),
            .I(N__36134));
    InMux I__6783 (
            .O(N__36200),
            .I(N__36134));
    InMux I__6782 (
            .O(N__36199),
            .I(N__36134));
    InMux I__6781 (
            .O(N__36198),
            .I(N__36134));
    InMux I__6780 (
            .O(N__36197),
            .I(N__36134));
    InMux I__6779 (
            .O(N__36196),
            .I(N__36125));
    InMux I__6778 (
            .O(N__36195),
            .I(N__36125));
    InMux I__6777 (
            .O(N__36194),
            .I(N__36125));
    InMux I__6776 (
            .O(N__36193),
            .I(N__36125));
    LocalMux I__6775 (
            .O(N__36184),
            .I(N__36114));
    LocalMux I__6774 (
            .O(N__36175),
            .I(N__36114));
    Span4Mux_v I__6773 (
            .O(N__36172),
            .I(N__36114));
    LocalMux I__6772 (
            .O(N__36163),
            .I(N__36114));
    LocalMux I__6771 (
            .O(N__36154),
            .I(N__36114));
    LocalMux I__6770 (
            .O(N__36145),
            .I(N__36109));
    LocalMux I__6769 (
            .O(N__36134),
            .I(N__36109));
    LocalMux I__6768 (
            .O(N__36125),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    Odrv4 I__6767 (
            .O(N__36114),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    Odrv12 I__6766 (
            .O(N__36109),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    InMux I__6765 (
            .O(N__36102),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_30 ));
    InMux I__6764 (
            .O(N__36099),
            .I(N__36094));
    InMux I__6763 (
            .O(N__36098),
            .I(N__36089));
    InMux I__6762 (
            .O(N__36097),
            .I(N__36089));
    LocalMux I__6761 (
            .O(N__36094),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    LocalMux I__6760 (
            .O(N__36089),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    CEMux I__6759 (
            .O(N__36084),
            .I(N__36081));
    LocalMux I__6758 (
            .O(N__36081),
            .I(N__36078));
    Span4Mux_v I__6757 (
            .O(N__36078),
            .I(N__36073));
    CEMux I__6756 (
            .O(N__36077),
            .I(N__36070));
    CEMux I__6755 (
            .O(N__36076),
            .I(N__36067));
    Span4Mux_v I__6754 (
            .O(N__36073),
            .I(N__36062));
    LocalMux I__6753 (
            .O(N__36070),
            .I(N__36062));
    LocalMux I__6752 (
            .O(N__36067),
            .I(N__36059));
    Span4Mux_v I__6751 (
            .O(N__36062),
            .I(N__36055));
    Span12Mux_h I__6750 (
            .O(N__36059),
            .I(N__36052));
    CEMux I__6749 (
            .O(N__36058),
            .I(N__36049));
    Odrv4 I__6748 (
            .O(N__36055),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv12 I__6747 (
            .O(N__36052),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__6746 (
            .O(N__36049),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__6745 (
            .O(N__36042),
            .I(N__36036));
    InMux I__6744 (
            .O(N__36041),
            .I(N__36036));
    LocalMux I__6743 (
            .O(N__36036),
            .I(N__36033));
    Odrv4 I__6742 (
            .O(N__36033),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ));
    InMux I__6741 (
            .O(N__36030),
            .I(N__36026));
    InMux I__6740 (
            .O(N__36029),
            .I(N__36023));
    LocalMux I__6739 (
            .O(N__36026),
            .I(N__36020));
    LocalMux I__6738 (
            .O(N__36023),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ));
    Odrv4 I__6737 (
            .O(N__36020),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ));
    InMux I__6736 (
            .O(N__36015),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_16 ));
    InMux I__6735 (
            .O(N__36012),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_17 ));
    InMux I__6734 (
            .O(N__36009),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_18 ));
    InMux I__6733 (
            .O(N__36006),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_19 ));
    InMux I__6732 (
            .O(N__36003),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_20 ));
    InMux I__6731 (
            .O(N__36000),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_21 ));
    InMux I__6730 (
            .O(N__35997),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_22 ));
    InMux I__6729 (
            .O(N__35994),
            .I(bfn_13_10_0_));
    InMux I__6728 (
            .O(N__35991),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_24 ));
    InMux I__6727 (
            .O(N__35988),
            .I(bfn_13_8_0_));
    InMux I__6726 (
            .O(N__35985),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_8 ));
    InMux I__6725 (
            .O(N__35982),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_9 ));
    InMux I__6724 (
            .O(N__35979),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_10 ));
    InMux I__6723 (
            .O(N__35976),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_11 ));
    InMux I__6722 (
            .O(N__35973),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_12 ));
    InMux I__6721 (
            .O(N__35970),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_13 ));
    InMux I__6720 (
            .O(N__35967),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_14 ));
    InMux I__6719 (
            .O(N__35964),
            .I(bfn_13_9_0_));
    InMux I__6718 (
            .O(N__35961),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_0 ));
    InMux I__6717 (
            .O(N__35958),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_1 ));
    InMux I__6716 (
            .O(N__35955),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_2 ));
    InMux I__6715 (
            .O(N__35952),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_3 ));
    InMux I__6714 (
            .O(N__35949),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_4 ));
    InMux I__6713 (
            .O(N__35946),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_5 ));
    InMux I__6712 (
            .O(N__35943),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_6 ));
    InMux I__6711 (
            .O(N__35940),
            .I(N__35935));
    InMux I__6710 (
            .O(N__35939),
            .I(N__35930));
    InMux I__6709 (
            .O(N__35938),
            .I(N__35930));
    LocalMux I__6708 (
            .O(N__35935),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    LocalMux I__6707 (
            .O(N__35930),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    InMux I__6706 (
            .O(N__35925),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_22 ));
    InMux I__6705 (
            .O(N__35922),
            .I(N__35917));
    InMux I__6704 (
            .O(N__35921),
            .I(N__35914));
    InMux I__6703 (
            .O(N__35920),
            .I(N__35911));
    LocalMux I__6702 (
            .O(N__35917),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    LocalMux I__6701 (
            .O(N__35914),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    LocalMux I__6700 (
            .O(N__35911),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    InMux I__6699 (
            .O(N__35904),
            .I(bfn_12_30_0_));
    CascadeMux I__6698 (
            .O(N__35901),
            .I(N__35897));
    InMux I__6697 (
            .O(N__35900),
            .I(N__35893));
    InMux I__6696 (
            .O(N__35897),
            .I(N__35890));
    InMux I__6695 (
            .O(N__35896),
            .I(N__35887));
    LocalMux I__6694 (
            .O(N__35893),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    LocalMux I__6693 (
            .O(N__35890),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    LocalMux I__6692 (
            .O(N__35887),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    InMux I__6691 (
            .O(N__35880),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_24 ));
    CascadeMux I__6690 (
            .O(N__35877),
            .I(N__35873));
    CascadeMux I__6689 (
            .O(N__35876),
            .I(N__35870));
    InMux I__6688 (
            .O(N__35873),
            .I(N__35867));
    InMux I__6687 (
            .O(N__35870),
            .I(N__35864));
    LocalMux I__6686 (
            .O(N__35867),
            .I(N__35858));
    LocalMux I__6685 (
            .O(N__35864),
            .I(N__35858));
    InMux I__6684 (
            .O(N__35863),
            .I(N__35855));
    Span4Mux_v I__6683 (
            .O(N__35858),
            .I(N__35852));
    LocalMux I__6682 (
            .O(N__35855),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ));
    Odrv4 I__6681 (
            .O(N__35852),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ));
    InMux I__6680 (
            .O(N__35847),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_25 ));
    InMux I__6679 (
            .O(N__35844),
            .I(N__35841));
    LocalMux I__6678 (
            .O(N__35841),
            .I(N__35836));
    InMux I__6677 (
            .O(N__35840),
            .I(N__35833));
    InMux I__6676 (
            .O(N__35839),
            .I(N__35830));
    Span4Mux_v I__6675 (
            .O(N__35836),
            .I(N__35827));
    LocalMux I__6674 (
            .O(N__35833),
            .I(N__35824));
    LocalMux I__6673 (
            .O(N__35830),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    Odrv4 I__6672 (
            .O(N__35827),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    Odrv12 I__6671 (
            .O(N__35824),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    InMux I__6670 (
            .O(N__35817),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_26 ));
    InMux I__6669 (
            .O(N__35814),
            .I(N__35810));
    InMux I__6668 (
            .O(N__35813),
            .I(N__35807));
    LocalMux I__6667 (
            .O(N__35810),
            .I(N__35801));
    LocalMux I__6666 (
            .O(N__35807),
            .I(N__35801));
    InMux I__6665 (
            .O(N__35806),
            .I(N__35798));
    Span4Mux_h I__6664 (
            .O(N__35801),
            .I(N__35795));
    LocalMux I__6663 (
            .O(N__35798),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ));
    Odrv4 I__6662 (
            .O(N__35795),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ));
    InMux I__6661 (
            .O(N__35790),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_27 ));
    InMux I__6660 (
            .O(N__35787),
            .I(N__35783));
    InMux I__6659 (
            .O(N__35786),
            .I(N__35779));
    LocalMux I__6658 (
            .O(N__35783),
            .I(N__35776));
    InMux I__6657 (
            .O(N__35782),
            .I(N__35773));
    LocalMux I__6656 (
            .O(N__35779),
            .I(N__35770));
    Span4Mux_h I__6655 (
            .O(N__35776),
            .I(N__35767));
    LocalMux I__6654 (
            .O(N__35773),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    Odrv4 I__6653 (
            .O(N__35770),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    Odrv4 I__6652 (
            .O(N__35767),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    InMux I__6651 (
            .O(N__35760),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_28 ));
    InMux I__6650 (
            .O(N__35757),
            .I(N__35752));
    InMux I__6649 (
            .O(N__35756),
            .I(N__35749));
    InMux I__6648 (
            .O(N__35755),
            .I(N__35746));
    LocalMux I__6647 (
            .O(N__35752),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    LocalMux I__6646 (
            .O(N__35749),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    LocalMux I__6645 (
            .O(N__35746),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    InMux I__6644 (
            .O(N__35739),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_29 ));
    InMux I__6643 (
            .O(N__35736),
            .I(N__35696));
    InMux I__6642 (
            .O(N__35735),
            .I(N__35696));
    InMux I__6641 (
            .O(N__35734),
            .I(N__35696));
    InMux I__6640 (
            .O(N__35733),
            .I(N__35696));
    InMux I__6639 (
            .O(N__35732),
            .I(N__35689));
    InMux I__6638 (
            .O(N__35731),
            .I(N__35689));
    InMux I__6637 (
            .O(N__35730),
            .I(N__35689));
    InMux I__6636 (
            .O(N__35729),
            .I(N__35680));
    InMux I__6635 (
            .O(N__35728),
            .I(N__35680));
    InMux I__6634 (
            .O(N__35727),
            .I(N__35680));
    InMux I__6633 (
            .O(N__35726),
            .I(N__35680));
    InMux I__6632 (
            .O(N__35725),
            .I(N__35669));
    InMux I__6631 (
            .O(N__35724),
            .I(N__35669));
    InMux I__6630 (
            .O(N__35723),
            .I(N__35669));
    InMux I__6629 (
            .O(N__35722),
            .I(N__35669));
    InMux I__6628 (
            .O(N__35721),
            .I(N__35669));
    InMux I__6627 (
            .O(N__35720),
            .I(N__35660));
    InMux I__6626 (
            .O(N__35719),
            .I(N__35660));
    InMux I__6625 (
            .O(N__35718),
            .I(N__35660));
    InMux I__6624 (
            .O(N__35717),
            .I(N__35660));
    InMux I__6623 (
            .O(N__35716),
            .I(N__35651));
    InMux I__6622 (
            .O(N__35715),
            .I(N__35651));
    InMux I__6621 (
            .O(N__35714),
            .I(N__35651));
    InMux I__6620 (
            .O(N__35713),
            .I(N__35651));
    InMux I__6619 (
            .O(N__35712),
            .I(N__35642));
    InMux I__6618 (
            .O(N__35711),
            .I(N__35642));
    InMux I__6617 (
            .O(N__35710),
            .I(N__35642));
    InMux I__6616 (
            .O(N__35709),
            .I(N__35642));
    InMux I__6615 (
            .O(N__35708),
            .I(N__35633));
    InMux I__6614 (
            .O(N__35707),
            .I(N__35633));
    InMux I__6613 (
            .O(N__35706),
            .I(N__35633));
    InMux I__6612 (
            .O(N__35705),
            .I(N__35633));
    LocalMux I__6611 (
            .O(N__35696),
            .I(N__35630));
    LocalMux I__6610 (
            .O(N__35689),
            .I(N__35627));
    LocalMux I__6609 (
            .O(N__35680),
            .I(N__35616));
    LocalMux I__6608 (
            .O(N__35669),
            .I(N__35616));
    LocalMux I__6607 (
            .O(N__35660),
            .I(N__35616));
    LocalMux I__6606 (
            .O(N__35651),
            .I(N__35616));
    LocalMux I__6605 (
            .O(N__35642),
            .I(N__35616));
    LocalMux I__6604 (
            .O(N__35633),
            .I(N__35613));
    Span4Mux_h I__6603 (
            .O(N__35630),
            .I(N__35606));
    Span4Mux_s3_v I__6602 (
            .O(N__35627),
            .I(N__35606));
    Span4Mux_s3_v I__6601 (
            .O(N__35616),
            .I(N__35606));
    Odrv12 I__6600 (
            .O(N__35613),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    Odrv4 I__6599 (
            .O(N__35606),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    InMux I__6598 (
            .O(N__35601),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_30 ));
    InMux I__6597 (
            .O(N__35598),
            .I(N__35593));
    InMux I__6596 (
            .O(N__35597),
            .I(N__35590));
    InMux I__6595 (
            .O(N__35596),
            .I(N__35587));
    LocalMux I__6594 (
            .O(N__35593),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    LocalMux I__6593 (
            .O(N__35590),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    LocalMux I__6592 (
            .O(N__35587),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    CEMux I__6591 (
            .O(N__35580),
            .I(N__35568));
    CEMux I__6590 (
            .O(N__35579),
            .I(N__35568));
    CEMux I__6589 (
            .O(N__35578),
            .I(N__35568));
    CEMux I__6588 (
            .O(N__35577),
            .I(N__35568));
    GlobalMux I__6587 (
            .O(N__35568),
            .I(N__35565));
    gio2CtrlBuf I__6586 (
            .O(N__35565),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_g ));
    InMux I__6585 (
            .O(N__35562),
            .I(N__35558));
    InMux I__6584 (
            .O(N__35561),
            .I(N__35555));
    LocalMux I__6583 (
            .O(N__35558),
            .I(N__35552));
    LocalMux I__6582 (
            .O(N__35555),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ));
    Odrv4 I__6581 (
            .O(N__35552),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ));
    InMux I__6580 (
            .O(N__35547),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_14 ));
    InMux I__6579 (
            .O(N__35544),
            .I(bfn_12_29_0_));
    InMux I__6578 (
            .O(N__35541),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_16 ));
    InMux I__6577 (
            .O(N__35538),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_17 ));
    InMux I__6576 (
            .O(N__35535),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_18 ));
    InMux I__6575 (
            .O(N__35532),
            .I(N__35527));
    InMux I__6574 (
            .O(N__35531),
            .I(N__35524));
    InMux I__6573 (
            .O(N__35530),
            .I(N__35521));
    LocalMux I__6572 (
            .O(N__35527),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    LocalMux I__6571 (
            .O(N__35524),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    LocalMux I__6570 (
            .O(N__35521),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    InMux I__6569 (
            .O(N__35514),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_19 ));
    CascadeMux I__6568 (
            .O(N__35511),
            .I(N__35507));
    InMux I__6567 (
            .O(N__35510),
            .I(N__35503));
    InMux I__6566 (
            .O(N__35507),
            .I(N__35500));
    InMux I__6565 (
            .O(N__35506),
            .I(N__35497));
    LocalMux I__6564 (
            .O(N__35503),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    LocalMux I__6563 (
            .O(N__35500),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    LocalMux I__6562 (
            .O(N__35497),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    InMux I__6561 (
            .O(N__35490),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_20 ));
    InMux I__6560 (
            .O(N__35487),
            .I(N__35482));
    InMux I__6559 (
            .O(N__35486),
            .I(N__35477));
    InMux I__6558 (
            .O(N__35485),
            .I(N__35477));
    LocalMux I__6557 (
            .O(N__35482),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    LocalMux I__6556 (
            .O(N__35477),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    InMux I__6555 (
            .O(N__35472),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_21 ));
    InMux I__6554 (
            .O(N__35469),
            .I(N__35465));
    InMux I__6553 (
            .O(N__35468),
            .I(N__35462));
    LocalMux I__6552 (
            .O(N__35465),
            .I(N__35459));
    LocalMux I__6551 (
            .O(N__35462),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ));
    Odrv4 I__6550 (
            .O(N__35459),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ));
    InMux I__6549 (
            .O(N__35454),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_5 ));
    InMux I__6548 (
            .O(N__35451),
            .I(N__35447));
    InMux I__6547 (
            .O(N__35450),
            .I(N__35444));
    LocalMux I__6546 (
            .O(N__35447),
            .I(N__35441));
    LocalMux I__6545 (
            .O(N__35444),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ));
    Odrv4 I__6544 (
            .O(N__35441),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ));
    InMux I__6543 (
            .O(N__35436),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_6 ));
    InMux I__6542 (
            .O(N__35433),
            .I(N__35429));
    InMux I__6541 (
            .O(N__35432),
            .I(N__35426));
    LocalMux I__6540 (
            .O(N__35429),
            .I(N__35423));
    LocalMux I__6539 (
            .O(N__35426),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ));
    Odrv4 I__6538 (
            .O(N__35423),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ));
    InMux I__6537 (
            .O(N__35418),
            .I(bfn_12_28_0_));
    InMux I__6536 (
            .O(N__35415),
            .I(N__35411));
    InMux I__6535 (
            .O(N__35414),
            .I(N__35408));
    LocalMux I__6534 (
            .O(N__35411),
            .I(N__35405));
    LocalMux I__6533 (
            .O(N__35408),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ));
    Odrv4 I__6532 (
            .O(N__35405),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ));
    InMux I__6531 (
            .O(N__35400),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_8 ));
    InMux I__6530 (
            .O(N__35397),
            .I(N__35393));
    InMux I__6529 (
            .O(N__35396),
            .I(N__35390));
    LocalMux I__6528 (
            .O(N__35393),
            .I(N__35387));
    LocalMux I__6527 (
            .O(N__35390),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ));
    Odrv4 I__6526 (
            .O(N__35387),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ));
    InMux I__6525 (
            .O(N__35382),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_9 ));
    InMux I__6524 (
            .O(N__35379),
            .I(N__35375));
    InMux I__6523 (
            .O(N__35378),
            .I(N__35372));
    LocalMux I__6522 (
            .O(N__35375),
            .I(N__35369));
    LocalMux I__6521 (
            .O(N__35372),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ));
    Odrv4 I__6520 (
            .O(N__35369),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ));
    InMux I__6519 (
            .O(N__35364),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_10 ));
    InMux I__6518 (
            .O(N__35361),
            .I(N__35357));
    InMux I__6517 (
            .O(N__35360),
            .I(N__35354));
    LocalMux I__6516 (
            .O(N__35357),
            .I(N__35351));
    LocalMux I__6515 (
            .O(N__35354),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ));
    Odrv4 I__6514 (
            .O(N__35351),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ));
    InMux I__6513 (
            .O(N__35346),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_11 ));
    InMux I__6512 (
            .O(N__35343),
            .I(N__35339));
    InMux I__6511 (
            .O(N__35342),
            .I(N__35336));
    LocalMux I__6510 (
            .O(N__35339),
            .I(N__35333));
    LocalMux I__6509 (
            .O(N__35336),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ));
    Odrv4 I__6508 (
            .O(N__35333),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ));
    InMux I__6507 (
            .O(N__35328),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_12 ));
    InMux I__6506 (
            .O(N__35325),
            .I(N__35321));
    InMux I__6505 (
            .O(N__35324),
            .I(N__35318));
    LocalMux I__6504 (
            .O(N__35321),
            .I(N__35315));
    LocalMux I__6503 (
            .O(N__35318),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ));
    Odrv4 I__6502 (
            .O(N__35315),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ));
    InMux I__6501 (
            .O(N__35310),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_13 ));
    InMux I__6500 (
            .O(N__35307),
            .I(N__35304));
    LocalMux I__6499 (
            .O(N__35304),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ));
    InMux I__6498 (
            .O(N__35301),
            .I(N__35297));
    InMux I__6497 (
            .O(N__35300),
            .I(N__35294));
    LocalMux I__6496 (
            .O(N__35297),
            .I(N__35291));
    LocalMux I__6495 (
            .O(N__35294),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ));
    Odrv4 I__6494 (
            .O(N__35291),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ));
    InMux I__6493 (
            .O(N__35286),
            .I(N__35282));
    InMux I__6492 (
            .O(N__35285),
            .I(N__35279));
    LocalMux I__6491 (
            .O(N__35282),
            .I(N__35276));
    LocalMux I__6490 (
            .O(N__35279),
            .I(N__35273));
    Odrv4 I__6489 (
            .O(N__35276),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ));
    Odrv12 I__6488 (
            .O(N__35273),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ));
    InMux I__6487 (
            .O(N__35268),
            .I(N__35265));
    LocalMux I__6486 (
            .O(N__35265),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__6485 (
            .O(N__35262),
            .I(N__35258));
    InMux I__6484 (
            .O(N__35261),
            .I(N__35255));
    InMux I__6483 (
            .O(N__35258),
            .I(N__35252));
    LocalMux I__6482 (
            .O(N__35255),
            .I(\phase_controller_inst1.stoper_tr.counter ));
    LocalMux I__6481 (
            .O(N__35252),
            .I(\phase_controller_inst1.stoper_tr.counter ));
    InMux I__6480 (
            .O(N__35247),
            .I(N__35243));
    InMux I__6479 (
            .O(N__35246),
            .I(N__35240));
    LocalMux I__6478 (
            .O(N__35243),
            .I(N__35237));
    LocalMux I__6477 (
            .O(N__35240),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ));
    Odrv4 I__6476 (
            .O(N__35237),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ));
    InMux I__6475 (
            .O(N__35232),
            .I(N__35228));
    InMux I__6474 (
            .O(N__35231),
            .I(N__35225));
    LocalMux I__6473 (
            .O(N__35228),
            .I(N__35222));
    LocalMux I__6472 (
            .O(N__35225),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ));
    Odrv4 I__6471 (
            .O(N__35222),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ));
    InMux I__6470 (
            .O(N__35217),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_0 ));
    InMux I__6469 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__6468 (
            .O(N__35211),
            .I(N__35207));
    InMux I__6467 (
            .O(N__35210),
            .I(N__35204));
    Span12Mux_h I__6466 (
            .O(N__35207),
            .I(N__35201));
    LocalMux I__6465 (
            .O(N__35204),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ));
    Odrv12 I__6464 (
            .O(N__35201),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ));
    InMux I__6463 (
            .O(N__35196),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_1 ));
    InMux I__6462 (
            .O(N__35193),
            .I(N__35190));
    LocalMux I__6461 (
            .O(N__35190),
            .I(N__35186));
    InMux I__6460 (
            .O(N__35189),
            .I(N__35183));
    Span4Mux_v I__6459 (
            .O(N__35186),
            .I(N__35180));
    LocalMux I__6458 (
            .O(N__35183),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ));
    Odrv4 I__6457 (
            .O(N__35180),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ));
    InMux I__6456 (
            .O(N__35175),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_2 ));
    InMux I__6455 (
            .O(N__35172),
            .I(N__35168));
    InMux I__6454 (
            .O(N__35171),
            .I(N__35165));
    LocalMux I__6453 (
            .O(N__35168),
            .I(N__35162));
    LocalMux I__6452 (
            .O(N__35165),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ));
    Odrv4 I__6451 (
            .O(N__35162),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ));
    InMux I__6450 (
            .O(N__35157),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_3 ));
    InMux I__6449 (
            .O(N__35154),
            .I(N__35151));
    LocalMux I__6448 (
            .O(N__35151),
            .I(N__35147));
    InMux I__6447 (
            .O(N__35150),
            .I(N__35144));
    Span4Mux_h I__6446 (
            .O(N__35147),
            .I(N__35141));
    LocalMux I__6445 (
            .O(N__35144),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ));
    Odrv4 I__6444 (
            .O(N__35141),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ));
    InMux I__6443 (
            .O(N__35136),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_4 ));
    InMux I__6442 (
            .O(N__35133),
            .I(N__35129));
    InMux I__6441 (
            .O(N__35132),
            .I(N__35126));
    LocalMux I__6440 (
            .O(N__35129),
            .I(N__35121));
    LocalMux I__6439 (
            .O(N__35126),
            .I(N__35121));
    Span4Mux_v I__6438 (
            .O(N__35121),
            .I(N__35118));
    Odrv4 I__6437 (
            .O(N__35118),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ));
    CascadeMux I__6436 (
            .O(N__35115),
            .I(N__35111));
    InMux I__6435 (
            .O(N__35114),
            .I(N__35108));
    InMux I__6434 (
            .O(N__35111),
            .I(N__35105));
    LocalMux I__6433 (
            .O(N__35108),
            .I(N__35100));
    LocalMux I__6432 (
            .O(N__35105),
            .I(N__35100));
    Span4Mux_v I__6431 (
            .O(N__35100),
            .I(N__35097));
    Odrv4 I__6430 (
            .O(N__35097),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ));
    InMux I__6429 (
            .O(N__35094),
            .I(N__35091));
    LocalMux I__6428 (
            .O(N__35091),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ));
    InMux I__6427 (
            .O(N__35088),
            .I(N__35085));
    LocalMux I__6426 (
            .O(N__35085),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ));
    InMux I__6425 (
            .O(N__35082),
            .I(N__35079));
    LocalMux I__6424 (
            .O(N__35079),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ));
    InMux I__6423 (
            .O(N__35076),
            .I(N__35073));
    LocalMux I__6422 (
            .O(N__35073),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ));
    InMux I__6421 (
            .O(N__35070),
            .I(N__35067));
    LocalMux I__6420 (
            .O(N__35067),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ));
    InMux I__6419 (
            .O(N__35064),
            .I(N__35061));
    LocalMux I__6418 (
            .O(N__35061),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ));
    InMux I__6417 (
            .O(N__35058),
            .I(N__35055));
    LocalMux I__6416 (
            .O(N__35055),
            .I(N__35052));
    Span4Mux_v I__6415 (
            .O(N__35052),
            .I(N__35049));
    Span4Mux_v I__6414 (
            .O(N__35049),
            .I(N__35046));
    Odrv4 I__6413 (
            .O(N__35046),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ));
    CascadeMux I__6412 (
            .O(N__35043),
            .I(N__35039));
    CascadeMux I__6411 (
            .O(N__35042),
            .I(N__35036));
    InMux I__6410 (
            .O(N__35039),
            .I(N__35031));
    InMux I__6409 (
            .O(N__35036),
            .I(N__35031));
    LocalMux I__6408 (
            .O(N__35031),
            .I(N__35028));
    Span4Mux_v I__6407 (
            .O(N__35028),
            .I(N__35025));
    Span4Mux_h I__6406 (
            .O(N__35025),
            .I(N__35022));
    Odrv4 I__6405 (
            .O(N__35022),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ));
    InMux I__6404 (
            .O(N__35019),
            .I(N__35016));
    LocalMux I__6403 (
            .O(N__35016),
            .I(N__35013));
    Span4Mux_v I__6402 (
            .O(N__35013),
            .I(N__35010));
    Odrv4 I__6401 (
            .O(N__35010),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ));
    InMux I__6400 (
            .O(N__35007),
            .I(N__35003));
    InMux I__6399 (
            .O(N__35006),
            .I(N__35000));
    LocalMux I__6398 (
            .O(N__35003),
            .I(N__34997));
    LocalMux I__6397 (
            .O(N__35000),
            .I(N__34994));
    Span4Mux_v I__6396 (
            .O(N__34997),
            .I(N__34989));
    Span4Mux_v I__6395 (
            .O(N__34994),
            .I(N__34989));
    Odrv4 I__6394 (
            .O(N__34989),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ));
    CascadeMux I__6393 (
            .O(N__34986),
            .I(N__34983));
    InMux I__6392 (
            .O(N__34983),
            .I(N__34980));
    LocalMux I__6391 (
            .O(N__34980),
            .I(N__34977));
    Span4Mux_v I__6390 (
            .O(N__34977),
            .I(N__34974));
    Odrv4 I__6389 (
            .O(N__34974),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ));
    CascadeMux I__6388 (
            .O(N__34971),
            .I(N__34967));
    InMux I__6387 (
            .O(N__34970),
            .I(N__34964));
    InMux I__6386 (
            .O(N__34967),
            .I(N__34961));
    LocalMux I__6385 (
            .O(N__34964),
            .I(N__34956));
    LocalMux I__6384 (
            .O(N__34961),
            .I(N__34956));
    Span4Mux_v I__6383 (
            .O(N__34956),
            .I(N__34953));
    Odrv4 I__6382 (
            .O(N__34953),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ));
    InMux I__6381 (
            .O(N__34950),
            .I(N__34946));
    CascadeMux I__6380 (
            .O(N__34949),
            .I(N__34941));
    LocalMux I__6379 (
            .O(N__34946),
            .I(N__34938));
    InMux I__6378 (
            .O(N__34945),
            .I(N__34935));
    InMux I__6377 (
            .O(N__34944),
            .I(N__34932));
    InMux I__6376 (
            .O(N__34941),
            .I(N__34929));
    Span4Mux_h I__6375 (
            .O(N__34938),
            .I(N__34926));
    LocalMux I__6374 (
            .O(N__34935),
            .I(N__34919));
    LocalMux I__6373 (
            .O(N__34932),
            .I(N__34919));
    LocalMux I__6372 (
            .O(N__34929),
            .I(N__34919));
    Span4Mux_v I__6371 (
            .O(N__34926),
            .I(N__34916));
    Span4Mux_v I__6370 (
            .O(N__34919),
            .I(N__34913));
    Odrv4 I__6369 (
            .O(N__34916),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ));
    Odrv4 I__6368 (
            .O(N__34913),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ));
    CascadeMux I__6367 (
            .O(N__34908),
            .I(N__34894));
    InMux I__6366 (
            .O(N__34907),
            .I(N__34888));
    InMux I__6365 (
            .O(N__34906),
            .I(N__34888));
    CascadeMux I__6364 (
            .O(N__34905),
            .I(N__34884));
    InMux I__6363 (
            .O(N__34904),
            .I(N__34871));
    InMux I__6362 (
            .O(N__34903),
            .I(N__34871));
    InMux I__6361 (
            .O(N__34902),
            .I(N__34871));
    InMux I__6360 (
            .O(N__34901),
            .I(N__34871));
    InMux I__6359 (
            .O(N__34900),
            .I(N__34871));
    InMux I__6358 (
            .O(N__34899),
            .I(N__34871));
    InMux I__6357 (
            .O(N__34898),
            .I(N__34866));
    InMux I__6356 (
            .O(N__34897),
            .I(N__34866));
    InMux I__6355 (
            .O(N__34894),
            .I(N__34861));
    InMux I__6354 (
            .O(N__34893),
            .I(N__34861));
    LocalMux I__6353 (
            .O(N__34888),
            .I(N__34840));
    InMux I__6352 (
            .O(N__34887),
            .I(N__34835));
    InMux I__6351 (
            .O(N__34884),
            .I(N__34835));
    LocalMux I__6350 (
            .O(N__34871),
            .I(N__34832));
    LocalMux I__6349 (
            .O(N__34866),
            .I(N__34827));
    LocalMux I__6348 (
            .O(N__34861),
            .I(N__34827));
    CascadeMux I__6347 (
            .O(N__34860),
            .I(N__34824));
    CascadeMux I__6346 (
            .O(N__34859),
            .I(N__34821));
    InMux I__6345 (
            .O(N__34858),
            .I(N__34818));
    InMux I__6344 (
            .O(N__34857),
            .I(N__34811));
    InMux I__6343 (
            .O(N__34856),
            .I(N__34811));
    InMux I__6342 (
            .O(N__34855),
            .I(N__34811));
    CascadeMux I__6341 (
            .O(N__34854),
            .I(N__34804));
    CascadeMux I__6340 (
            .O(N__34853),
            .I(N__34801));
    CascadeMux I__6339 (
            .O(N__34852),
            .I(N__34794));
    CascadeMux I__6338 (
            .O(N__34851),
            .I(N__34788));
    CascadeMux I__6337 (
            .O(N__34850),
            .I(N__34779));
    CascadeMux I__6336 (
            .O(N__34849),
            .I(N__34776));
    CascadeMux I__6335 (
            .O(N__34848),
            .I(N__34769));
    CascadeMux I__6334 (
            .O(N__34847),
            .I(N__34766));
    CascadeMux I__6333 (
            .O(N__34846),
            .I(N__34759));
    CascadeMux I__6332 (
            .O(N__34845),
            .I(N__34755));
    CascadeMux I__6331 (
            .O(N__34844),
            .I(N__34751));
    CascadeMux I__6330 (
            .O(N__34843),
            .I(N__34747));
    Span4Mux_h I__6329 (
            .O(N__34840),
            .I(N__34726));
    LocalMux I__6328 (
            .O(N__34835),
            .I(N__34726));
    Span4Mux_h I__6327 (
            .O(N__34832),
            .I(N__34726));
    Span4Mux_v I__6326 (
            .O(N__34827),
            .I(N__34723));
    InMux I__6325 (
            .O(N__34824),
            .I(N__34720));
    InMux I__6324 (
            .O(N__34821),
            .I(N__34717));
    LocalMux I__6323 (
            .O(N__34818),
            .I(N__34712));
    LocalMux I__6322 (
            .O(N__34811),
            .I(N__34712));
    InMux I__6321 (
            .O(N__34810),
            .I(N__34703));
    InMux I__6320 (
            .O(N__34809),
            .I(N__34703));
    InMux I__6319 (
            .O(N__34808),
            .I(N__34703));
    InMux I__6318 (
            .O(N__34807),
            .I(N__34703));
    InMux I__6317 (
            .O(N__34804),
            .I(N__34700));
    InMux I__6316 (
            .O(N__34801),
            .I(N__34697));
    InMux I__6315 (
            .O(N__34800),
            .I(N__34686));
    InMux I__6314 (
            .O(N__34799),
            .I(N__34686));
    InMux I__6313 (
            .O(N__34798),
            .I(N__34686));
    InMux I__6312 (
            .O(N__34797),
            .I(N__34686));
    InMux I__6311 (
            .O(N__34794),
            .I(N__34686));
    CascadeMux I__6310 (
            .O(N__34793),
            .I(N__34678));
    CascadeMux I__6309 (
            .O(N__34792),
            .I(N__34673));
    CascadeMux I__6308 (
            .O(N__34791),
            .I(N__34670));
    InMux I__6307 (
            .O(N__34788),
            .I(N__34667));
    InMux I__6306 (
            .O(N__34787),
            .I(N__34664));
    CascadeMux I__6305 (
            .O(N__34786),
            .I(N__34661));
    CascadeMux I__6304 (
            .O(N__34785),
            .I(N__34658));
    InMux I__6303 (
            .O(N__34784),
            .I(N__34647));
    InMux I__6302 (
            .O(N__34783),
            .I(N__34647));
    InMux I__6301 (
            .O(N__34782),
            .I(N__34647));
    InMux I__6300 (
            .O(N__34779),
            .I(N__34647));
    InMux I__6299 (
            .O(N__34776),
            .I(N__34647));
    InMux I__6298 (
            .O(N__34775),
            .I(N__34644));
    InMux I__6297 (
            .O(N__34774),
            .I(N__34630));
    InMux I__6296 (
            .O(N__34773),
            .I(N__34630));
    InMux I__6295 (
            .O(N__34772),
            .I(N__34630));
    InMux I__6294 (
            .O(N__34769),
            .I(N__34625));
    InMux I__6293 (
            .O(N__34766),
            .I(N__34625));
    CascadeMux I__6292 (
            .O(N__34765),
            .I(N__34622));
    CascadeMux I__6291 (
            .O(N__34764),
            .I(N__34618));
    CascadeMux I__6290 (
            .O(N__34763),
            .I(N__34614));
    InMux I__6289 (
            .O(N__34762),
            .I(N__34596));
    InMux I__6288 (
            .O(N__34759),
            .I(N__34596));
    InMux I__6287 (
            .O(N__34758),
            .I(N__34596));
    InMux I__6286 (
            .O(N__34755),
            .I(N__34596));
    InMux I__6285 (
            .O(N__34754),
            .I(N__34596));
    InMux I__6284 (
            .O(N__34751),
            .I(N__34596));
    InMux I__6283 (
            .O(N__34750),
            .I(N__34596));
    InMux I__6282 (
            .O(N__34747),
            .I(N__34596));
    CascadeMux I__6281 (
            .O(N__34746),
            .I(N__34593));
    CascadeMux I__6280 (
            .O(N__34745),
            .I(N__34589));
    CascadeMux I__6279 (
            .O(N__34744),
            .I(N__34585));
    CascadeMux I__6278 (
            .O(N__34743),
            .I(N__34581));
    CascadeMux I__6277 (
            .O(N__34742),
            .I(N__34577));
    CascadeMux I__6276 (
            .O(N__34741),
            .I(N__34573));
    CascadeMux I__6275 (
            .O(N__34740),
            .I(N__34569));
    CascadeMux I__6274 (
            .O(N__34739),
            .I(N__34565));
    CascadeMux I__6273 (
            .O(N__34738),
            .I(N__34560));
    CascadeMux I__6272 (
            .O(N__34737),
            .I(N__34556));
    CascadeMux I__6271 (
            .O(N__34736),
            .I(N__34552));
    CascadeMux I__6270 (
            .O(N__34735),
            .I(N__34547));
    CascadeMux I__6269 (
            .O(N__34734),
            .I(N__34543));
    CascadeMux I__6268 (
            .O(N__34733),
            .I(N__34539));
    Span4Mux_v I__6267 (
            .O(N__34726),
            .I(N__34529));
    Span4Mux_h I__6266 (
            .O(N__34723),
            .I(N__34529));
    LocalMux I__6265 (
            .O(N__34720),
            .I(N__34529));
    LocalMux I__6264 (
            .O(N__34717),
            .I(N__34529));
    Span4Mux_v I__6263 (
            .O(N__34712),
            .I(N__34526));
    LocalMux I__6262 (
            .O(N__34703),
            .I(N__34517));
    LocalMux I__6261 (
            .O(N__34700),
            .I(N__34517));
    LocalMux I__6260 (
            .O(N__34697),
            .I(N__34517));
    LocalMux I__6259 (
            .O(N__34686),
            .I(N__34517));
    InMux I__6258 (
            .O(N__34685),
            .I(N__34508));
    InMux I__6257 (
            .O(N__34684),
            .I(N__34508));
    InMux I__6256 (
            .O(N__34683),
            .I(N__34508));
    InMux I__6255 (
            .O(N__34682),
            .I(N__34508));
    InMux I__6254 (
            .O(N__34681),
            .I(N__34505));
    InMux I__6253 (
            .O(N__34678),
            .I(N__34494));
    InMux I__6252 (
            .O(N__34677),
            .I(N__34494));
    InMux I__6251 (
            .O(N__34676),
            .I(N__34494));
    InMux I__6250 (
            .O(N__34673),
            .I(N__34494));
    InMux I__6249 (
            .O(N__34670),
            .I(N__34494));
    LocalMux I__6248 (
            .O(N__34667),
            .I(N__34485));
    LocalMux I__6247 (
            .O(N__34664),
            .I(N__34485));
    InMux I__6246 (
            .O(N__34661),
            .I(N__34482));
    InMux I__6245 (
            .O(N__34658),
            .I(N__34479));
    LocalMux I__6244 (
            .O(N__34647),
            .I(N__34474));
    LocalMux I__6243 (
            .O(N__34644),
            .I(N__34474));
    CascadeMux I__6242 (
            .O(N__34643),
            .I(N__34471));
    CascadeMux I__6241 (
            .O(N__34642),
            .I(N__34467));
    CascadeMux I__6240 (
            .O(N__34641),
            .I(N__34463));
    CascadeMux I__6239 (
            .O(N__34640),
            .I(N__34459));
    CascadeMux I__6238 (
            .O(N__34639),
            .I(N__34455));
    CascadeMux I__6237 (
            .O(N__34638),
            .I(N__34451));
    CascadeMux I__6236 (
            .O(N__34637),
            .I(N__34447));
    LocalMux I__6235 (
            .O(N__34630),
            .I(N__34441));
    LocalMux I__6234 (
            .O(N__34625),
            .I(N__34441));
    InMux I__6233 (
            .O(N__34622),
            .I(N__34428));
    InMux I__6232 (
            .O(N__34621),
            .I(N__34428));
    InMux I__6231 (
            .O(N__34618),
            .I(N__34428));
    InMux I__6230 (
            .O(N__34617),
            .I(N__34428));
    InMux I__6229 (
            .O(N__34614),
            .I(N__34428));
    InMux I__6228 (
            .O(N__34613),
            .I(N__34428));
    LocalMux I__6227 (
            .O(N__34596),
            .I(N__34425));
    InMux I__6226 (
            .O(N__34593),
            .I(N__34408));
    InMux I__6225 (
            .O(N__34592),
            .I(N__34408));
    InMux I__6224 (
            .O(N__34589),
            .I(N__34408));
    InMux I__6223 (
            .O(N__34588),
            .I(N__34408));
    InMux I__6222 (
            .O(N__34585),
            .I(N__34408));
    InMux I__6221 (
            .O(N__34584),
            .I(N__34408));
    InMux I__6220 (
            .O(N__34581),
            .I(N__34408));
    InMux I__6219 (
            .O(N__34580),
            .I(N__34408));
    InMux I__6218 (
            .O(N__34577),
            .I(N__34391));
    InMux I__6217 (
            .O(N__34576),
            .I(N__34391));
    InMux I__6216 (
            .O(N__34573),
            .I(N__34391));
    InMux I__6215 (
            .O(N__34572),
            .I(N__34391));
    InMux I__6214 (
            .O(N__34569),
            .I(N__34391));
    InMux I__6213 (
            .O(N__34568),
            .I(N__34391));
    InMux I__6212 (
            .O(N__34565),
            .I(N__34391));
    InMux I__6211 (
            .O(N__34564),
            .I(N__34391));
    InMux I__6210 (
            .O(N__34563),
            .I(N__34376));
    InMux I__6209 (
            .O(N__34560),
            .I(N__34376));
    InMux I__6208 (
            .O(N__34559),
            .I(N__34376));
    InMux I__6207 (
            .O(N__34556),
            .I(N__34376));
    InMux I__6206 (
            .O(N__34555),
            .I(N__34376));
    InMux I__6205 (
            .O(N__34552),
            .I(N__34376));
    InMux I__6204 (
            .O(N__34551),
            .I(N__34376));
    InMux I__6203 (
            .O(N__34550),
            .I(N__34373));
    InMux I__6202 (
            .O(N__34547),
            .I(N__34360));
    InMux I__6201 (
            .O(N__34546),
            .I(N__34360));
    InMux I__6200 (
            .O(N__34543),
            .I(N__34360));
    InMux I__6199 (
            .O(N__34542),
            .I(N__34360));
    InMux I__6198 (
            .O(N__34539),
            .I(N__34360));
    InMux I__6197 (
            .O(N__34538),
            .I(N__34360));
    Span4Mux_v I__6196 (
            .O(N__34529),
            .I(N__34357));
    Span4Mux_h I__6195 (
            .O(N__34526),
            .I(N__34346));
    Span4Mux_v I__6194 (
            .O(N__34517),
            .I(N__34346));
    LocalMux I__6193 (
            .O(N__34508),
            .I(N__34346));
    LocalMux I__6192 (
            .O(N__34505),
            .I(N__34346));
    LocalMux I__6191 (
            .O(N__34494),
            .I(N__34346));
    InMux I__6190 (
            .O(N__34493),
            .I(N__34337));
    InMux I__6189 (
            .O(N__34492),
            .I(N__34337));
    InMux I__6188 (
            .O(N__34491),
            .I(N__34337));
    InMux I__6187 (
            .O(N__34490),
            .I(N__34337));
    Span4Mux_v I__6186 (
            .O(N__34485),
            .I(N__34328));
    LocalMux I__6185 (
            .O(N__34482),
            .I(N__34328));
    LocalMux I__6184 (
            .O(N__34479),
            .I(N__34328));
    Span4Mux_h I__6183 (
            .O(N__34474),
            .I(N__34328));
    InMux I__6182 (
            .O(N__34471),
            .I(N__34311));
    InMux I__6181 (
            .O(N__34470),
            .I(N__34311));
    InMux I__6180 (
            .O(N__34467),
            .I(N__34311));
    InMux I__6179 (
            .O(N__34466),
            .I(N__34311));
    InMux I__6178 (
            .O(N__34463),
            .I(N__34311));
    InMux I__6177 (
            .O(N__34462),
            .I(N__34311));
    InMux I__6176 (
            .O(N__34459),
            .I(N__34311));
    InMux I__6175 (
            .O(N__34458),
            .I(N__34311));
    InMux I__6174 (
            .O(N__34455),
            .I(N__34298));
    InMux I__6173 (
            .O(N__34454),
            .I(N__34298));
    InMux I__6172 (
            .O(N__34451),
            .I(N__34298));
    InMux I__6171 (
            .O(N__34450),
            .I(N__34298));
    InMux I__6170 (
            .O(N__34447),
            .I(N__34298));
    InMux I__6169 (
            .O(N__34446),
            .I(N__34298));
    Sp12to4 I__6168 (
            .O(N__34441),
            .I(N__34281));
    LocalMux I__6167 (
            .O(N__34428),
            .I(N__34281));
    Span12Mux_s9_v I__6166 (
            .O(N__34425),
            .I(N__34281));
    LocalMux I__6165 (
            .O(N__34408),
            .I(N__34281));
    LocalMux I__6164 (
            .O(N__34391),
            .I(N__34281));
    LocalMux I__6163 (
            .O(N__34376),
            .I(N__34281));
    LocalMux I__6162 (
            .O(N__34373),
            .I(N__34281));
    LocalMux I__6161 (
            .O(N__34360),
            .I(N__34281));
    Odrv4 I__6160 (
            .O(N__34357),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6159 (
            .O(N__34346),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6158 (
            .O(N__34337),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6157 (
            .O(N__34328),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6156 (
            .O(N__34311),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6155 (
            .O(N__34298),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__6154 (
            .O(N__34281),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__6153 (
            .O(N__34266),
            .I(N__34261));
    InMux I__6152 (
            .O(N__34265),
            .I(N__34255));
    InMux I__6151 (
            .O(N__34264),
            .I(N__34247));
    InMux I__6150 (
            .O(N__34261),
            .I(N__34247));
    InMux I__6149 (
            .O(N__34260),
            .I(N__34247));
    InMux I__6148 (
            .O(N__34259),
            .I(N__34239));
    InMux I__6147 (
            .O(N__34258),
            .I(N__34231));
    LocalMux I__6146 (
            .O(N__34255),
            .I(N__34226));
    InMux I__6145 (
            .O(N__34254),
            .I(N__34223));
    LocalMux I__6144 (
            .O(N__34247),
            .I(N__34220));
    InMux I__6143 (
            .O(N__34246),
            .I(N__34215));
    InMux I__6142 (
            .O(N__34245),
            .I(N__34215));
    InMux I__6141 (
            .O(N__34244),
            .I(N__34212));
    InMux I__6140 (
            .O(N__34243),
            .I(N__34203));
    InMux I__6139 (
            .O(N__34242),
            .I(N__34203));
    LocalMux I__6138 (
            .O(N__34239),
            .I(N__34182));
    InMux I__6137 (
            .O(N__34238),
            .I(N__34177));
    InMux I__6136 (
            .O(N__34237),
            .I(N__34177));
    InMux I__6135 (
            .O(N__34236),
            .I(N__34174));
    InMux I__6134 (
            .O(N__34235),
            .I(N__34169));
    InMux I__6133 (
            .O(N__34234),
            .I(N__34169));
    LocalMux I__6132 (
            .O(N__34231),
            .I(N__34166));
    InMux I__6131 (
            .O(N__34230),
            .I(N__34163));
    InMux I__6130 (
            .O(N__34229),
            .I(N__34160));
    Span4Mux_v I__6129 (
            .O(N__34226),
            .I(N__34153));
    LocalMux I__6128 (
            .O(N__34223),
            .I(N__34153));
    Span4Mux_h I__6127 (
            .O(N__34220),
            .I(N__34153));
    LocalMux I__6126 (
            .O(N__34215),
            .I(N__34148));
    LocalMux I__6125 (
            .O(N__34212),
            .I(N__34148));
    InMux I__6124 (
            .O(N__34211),
            .I(N__34141));
    InMux I__6123 (
            .O(N__34210),
            .I(N__34141));
    InMux I__6122 (
            .O(N__34209),
            .I(N__34141));
    InMux I__6121 (
            .O(N__34208),
            .I(N__34138));
    LocalMux I__6120 (
            .O(N__34203),
            .I(N__34130));
    InMux I__6119 (
            .O(N__34202),
            .I(N__34117));
    InMux I__6118 (
            .O(N__34201),
            .I(N__34117));
    InMux I__6117 (
            .O(N__34200),
            .I(N__34117));
    InMux I__6116 (
            .O(N__34199),
            .I(N__34117));
    InMux I__6115 (
            .O(N__34198),
            .I(N__34117));
    InMux I__6114 (
            .O(N__34197),
            .I(N__34117));
    InMux I__6113 (
            .O(N__34196),
            .I(N__34100));
    InMux I__6112 (
            .O(N__34195),
            .I(N__34100));
    InMux I__6111 (
            .O(N__34194),
            .I(N__34100));
    InMux I__6110 (
            .O(N__34193),
            .I(N__34100));
    InMux I__6109 (
            .O(N__34192),
            .I(N__34100));
    InMux I__6108 (
            .O(N__34191),
            .I(N__34100));
    InMux I__6107 (
            .O(N__34190),
            .I(N__34100));
    InMux I__6106 (
            .O(N__34189),
            .I(N__34100));
    InMux I__6105 (
            .O(N__34188),
            .I(N__34091));
    InMux I__6104 (
            .O(N__34187),
            .I(N__34091));
    InMux I__6103 (
            .O(N__34186),
            .I(N__34091));
    InMux I__6102 (
            .O(N__34185),
            .I(N__34091));
    Span4Mux_v I__6101 (
            .O(N__34182),
            .I(N__34083));
    LocalMux I__6100 (
            .O(N__34177),
            .I(N__34080));
    LocalMux I__6099 (
            .O(N__34174),
            .I(N__34057));
    LocalMux I__6098 (
            .O(N__34169),
            .I(N__34046));
    Span4Mux_h I__6097 (
            .O(N__34166),
            .I(N__34046));
    LocalMux I__6096 (
            .O(N__34163),
            .I(N__34046));
    LocalMux I__6095 (
            .O(N__34160),
            .I(N__34046));
    Span4Mux_v I__6094 (
            .O(N__34153),
            .I(N__34046));
    Span4Mux_v I__6093 (
            .O(N__34148),
            .I(N__34039));
    LocalMux I__6092 (
            .O(N__34141),
            .I(N__34039));
    LocalMux I__6091 (
            .O(N__34138),
            .I(N__34039));
    InMux I__6090 (
            .O(N__34137),
            .I(N__34034));
    InMux I__6089 (
            .O(N__34136),
            .I(N__34034));
    InMux I__6088 (
            .O(N__34135),
            .I(N__34027));
    InMux I__6087 (
            .O(N__34134),
            .I(N__34027));
    InMux I__6086 (
            .O(N__34133),
            .I(N__34027));
    Span4Mux_h I__6085 (
            .O(N__34130),
            .I(N__34018));
    LocalMux I__6084 (
            .O(N__34117),
            .I(N__34018));
    LocalMux I__6083 (
            .O(N__34100),
            .I(N__34018));
    LocalMux I__6082 (
            .O(N__34091),
            .I(N__34018));
    InMux I__6081 (
            .O(N__34090),
            .I(N__34015));
    InMux I__6080 (
            .O(N__34089),
            .I(N__34006));
    InMux I__6079 (
            .O(N__34088),
            .I(N__34006));
    InMux I__6078 (
            .O(N__34087),
            .I(N__34006));
    InMux I__6077 (
            .O(N__34086),
            .I(N__34006));
    Span4Mux_h I__6076 (
            .O(N__34083),
            .I(N__34001));
    Span4Mux_v I__6075 (
            .O(N__34080),
            .I(N__34001));
    InMux I__6074 (
            .O(N__34079),
            .I(N__33998));
    InMux I__6073 (
            .O(N__34078),
            .I(N__33985));
    InMux I__6072 (
            .O(N__34077),
            .I(N__33985));
    InMux I__6071 (
            .O(N__34076),
            .I(N__33985));
    InMux I__6070 (
            .O(N__34075),
            .I(N__33985));
    InMux I__6069 (
            .O(N__34074),
            .I(N__33985));
    InMux I__6068 (
            .O(N__34073),
            .I(N__33985));
    InMux I__6067 (
            .O(N__34072),
            .I(N__33974));
    InMux I__6066 (
            .O(N__34071),
            .I(N__33974));
    InMux I__6065 (
            .O(N__34070),
            .I(N__33974));
    InMux I__6064 (
            .O(N__34069),
            .I(N__33974));
    InMux I__6063 (
            .O(N__34068),
            .I(N__33974));
    InMux I__6062 (
            .O(N__34067),
            .I(N__33961));
    InMux I__6061 (
            .O(N__34066),
            .I(N__33961));
    InMux I__6060 (
            .O(N__34065),
            .I(N__33961));
    InMux I__6059 (
            .O(N__34064),
            .I(N__33961));
    InMux I__6058 (
            .O(N__34063),
            .I(N__33961));
    InMux I__6057 (
            .O(N__34062),
            .I(N__33961));
    InMux I__6056 (
            .O(N__34061),
            .I(N__33956));
    InMux I__6055 (
            .O(N__34060),
            .I(N__33956));
    Span4Mux_h I__6054 (
            .O(N__34057),
            .I(N__33949));
    Span4Mux_v I__6053 (
            .O(N__34046),
            .I(N__33949));
    Span4Mux_v I__6052 (
            .O(N__34039),
            .I(N__33949));
    LocalMux I__6051 (
            .O(N__34034),
            .I(N__33942));
    LocalMux I__6050 (
            .O(N__34027),
            .I(N__33942));
    Span4Mux_v I__6049 (
            .O(N__34018),
            .I(N__33942));
    LocalMux I__6048 (
            .O(N__34015),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6047 (
            .O(N__34006),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6046 (
            .O(N__34001),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6045 (
            .O(N__33998),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6044 (
            .O(N__33985),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6043 (
            .O(N__33974),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6042 (
            .O(N__33961),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6041 (
            .O(N__33956),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6040 (
            .O(N__33949),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6039 (
            .O(N__33942),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__6038 (
            .O(N__33921),
            .I(N__33918));
    InMux I__6037 (
            .O(N__33918),
            .I(N__33912));
    InMux I__6036 (
            .O(N__33917),
            .I(N__33907));
    InMux I__6035 (
            .O(N__33916),
            .I(N__33907));
    InMux I__6034 (
            .O(N__33915),
            .I(N__33904));
    LocalMux I__6033 (
            .O(N__33912),
            .I(N__33901));
    LocalMux I__6032 (
            .O(N__33907),
            .I(N__33898));
    LocalMux I__6031 (
            .O(N__33904),
            .I(N__33895));
    Span4Mux_v I__6030 (
            .O(N__33901),
            .I(N__33892));
    Span4Mux_v I__6029 (
            .O(N__33898),
            .I(N__33887));
    Span4Mux_h I__6028 (
            .O(N__33895),
            .I(N__33887));
    Odrv4 I__6027 (
            .O(N__33892),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__6026 (
            .O(N__33887),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__6025 (
            .O(N__33882),
            .I(N__33877));
    InMux I__6024 (
            .O(N__33881),
            .I(N__33872));
    InMux I__6023 (
            .O(N__33880),
            .I(N__33872));
    LocalMux I__6022 (
            .O(N__33877),
            .I(N__33869));
    LocalMux I__6021 (
            .O(N__33872),
            .I(N__33866));
    Odrv4 I__6020 (
            .O(N__33869),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__6019 (
            .O(N__33866),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__6018 (
            .O(N__33861),
            .I(N__33858));
    LocalMux I__6017 (
            .O(N__33858),
            .I(N__33855));
    Span4Mux_h I__6016 (
            .O(N__33855),
            .I(N__33852));
    Odrv4 I__6015 (
            .O(N__33852),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__6014 (
            .O(N__33849),
            .I(N__33846));
    LocalMux I__6013 (
            .O(N__33846),
            .I(N__33843));
    Sp12to4 I__6012 (
            .O(N__33843),
            .I(N__33840));
    Odrv12 I__6011 (
            .O(N__33840),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ));
    InMux I__6010 (
            .O(N__33837),
            .I(N__33834));
    LocalMux I__6009 (
            .O(N__33834),
            .I(N__33831));
    Span4Mux_v I__6008 (
            .O(N__33831),
            .I(N__33828));
    Odrv4 I__6007 (
            .O(N__33828),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ));
    InMux I__6006 (
            .O(N__33825),
            .I(N__33822));
    LocalMux I__6005 (
            .O(N__33822),
            .I(N__33819));
    Span4Mux_v I__6004 (
            .O(N__33819),
            .I(N__33816));
    Odrv4 I__6003 (
            .O(N__33816),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ));
    InMux I__6002 (
            .O(N__33813),
            .I(N__33810));
    LocalMux I__6001 (
            .O(N__33810),
            .I(N__33807));
    Span4Mux_v I__6000 (
            .O(N__33807),
            .I(N__33804));
    Odrv4 I__5999 (
            .O(N__33804),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ));
    InMux I__5998 (
            .O(N__33801),
            .I(N__33798));
    LocalMux I__5997 (
            .O(N__33798),
            .I(N__33795));
    Span4Mux_v I__5996 (
            .O(N__33795),
            .I(N__33792));
    Odrv4 I__5995 (
            .O(N__33792),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ));
    InMux I__5994 (
            .O(N__33789),
            .I(N__33786));
    LocalMux I__5993 (
            .O(N__33786),
            .I(N__33783));
    Span4Mux_v I__5992 (
            .O(N__33783),
            .I(N__33780));
    Odrv4 I__5991 (
            .O(N__33780),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ));
    InMux I__5990 (
            .O(N__33777),
            .I(N__33771));
    InMux I__5989 (
            .O(N__33776),
            .I(N__33771));
    LocalMux I__5988 (
            .O(N__33771),
            .I(N__33768));
    Span4Mux_h I__5987 (
            .O(N__33768),
            .I(N__33765));
    Span4Mux_v I__5986 (
            .O(N__33765),
            .I(N__33762));
    Odrv4 I__5985 (
            .O(N__33762),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ));
    CEMux I__5984 (
            .O(N__33759),
            .I(N__33735));
    CEMux I__5983 (
            .O(N__33758),
            .I(N__33735));
    CEMux I__5982 (
            .O(N__33757),
            .I(N__33735));
    CEMux I__5981 (
            .O(N__33756),
            .I(N__33735));
    CEMux I__5980 (
            .O(N__33755),
            .I(N__33735));
    CEMux I__5979 (
            .O(N__33754),
            .I(N__33735));
    CEMux I__5978 (
            .O(N__33753),
            .I(N__33735));
    CEMux I__5977 (
            .O(N__33752),
            .I(N__33735));
    GlobalMux I__5976 (
            .O(N__33735),
            .I(N__33732));
    gio2CtrlBuf I__5975 (
            .O(N__33732),
            .I(\current_shift_inst.timer_s1.N_153_i_g ));
    InMux I__5974 (
            .O(N__33729),
            .I(N__33726));
    LocalMux I__5973 (
            .O(N__33726),
            .I(N__33723));
    Span4Mux_v I__5972 (
            .O(N__33723),
            .I(N__33719));
    InMux I__5971 (
            .O(N__33722),
            .I(N__33716));
    Odrv4 I__5970 (
            .O(N__33719),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    LocalMux I__5969 (
            .O(N__33716),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__5968 (
            .O(N__33711),
            .I(N__33708));
    InMux I__5967 (
            .O(N__33708),
            .I(N__33705));
    LocalMux I__5966 (
            .O(N__33705),
            .I(N__33702));
    Span4Mux_v I__5965 (
            .O(N__33702),
            .I(N__33699));
    Odrv4 I__5964 (
            .O(N__33699),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__5963 (
            .O(N__33696),
            .I(N__33693));
    LocalMux I__5962 (
            .O(N__33693),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    CascadeMux I__5961 (
            .O(N__33690),
            .I(N__33686));
    CascadeMux I__5960 (
            .O(N__33689),
            .I(N__33683));
    InMux I__5959 (
            .O(N__33686),
            .I(N__33679));
    InMux I__5958 (
            .O(N__33683),
            .I(N__33676));
    InMux I__5957 (
            .O(N__33682),
            .I(N__33673));
    LocalMux I__5956 (
            .O(N__33679),
            .I(N__33670));
    LocalMux I__5955 (
            .O(N__33676),
            .I(N__33666));
    LocalMux I__5954 (
            .O(N__33673),
            .I(N__33663));
    Span4Mux_v I__5953 (
            .O(N__33670),
            .I(N__33660));
    InMux I__5952 (
            .O(N__33669),
            .I(N__33657));
    Span4Mux_h I__5951 (
            .O(N__33666),
            .I(N__33652));
    Span4Mux_v I__5950 (
            .O(N__33663),
            .I(N__33652));
    Sp12to4 I__5949 (
            .O(N__33660),
            .I(N__33647));
    LocalMux I__5948 (
            .O(N__33657),
            .I(N__33647));
    Odrv4 I__5947 (
            .O(N__33652),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv12 I__5946 (
            .O(N__33647),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__5945 (
            .O(N__33642),
            .I(N__33639));
    LocalMux I__5944 (
            .O(N__33639),
            .I(N__33634));
    InMux I__5943 (
            .O(N__33638),
            .I(N__33631));
    InMux I__5942 (
            .O(N__33637),
            .I(N__33628));
    Span4Mux_h I__5941 (
            .O(N__33634),
            .I(N__33625));
    LocalMux I__5940 (
            .O(N__33631),
            .I(N__33622));
    LocalMux I__5939 (
            .O(N__33628),
            .I(N__33619));
    Odrv4 I__5938 (
            .O(N__33625),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__5937 (
            .O(N__33622),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__5936 (
            .O(N__33619),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__5935 (
            .O(N__33612),
            .I(N__33609));
    LocalMux I__5934 (
            .O(N__33609),
            .I(N__33606));
    Span4Mux_h I__5933 (
            .O(N__33606),
            .I(N__33603));
    Odrv4 I__5932 (
            .O(N__33603),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    CascadeMux I__5931 (
            .O(N__33600),
            .I(N__33597));
    InMux I__5930 (
            .O(N__33597),
            .I(N__33593));
    CascadeMux I__5929 (
            .O(N__33596),
            .I(N__33590));
    LocalMux I__5928 (
            .O(N__33593),
            .I(N__33585));
    InMux I__5927 (
            .O(N__33590),
            .I(N__33582));
    InMux I__5926 (
            .O(N__33589),
            .I(N__33579));
    InMux I__5925 (
            .O(N__33588),
            .I(N__33576));
    Span4Mux_v I__5924 (
            .O(N__33585),
            .I(N__33569));
    LocalMux I__5923 (
            .O(N__33582),
            .I(N__33569));
    LocalMux I__5922 (
            .O(N__33579),
            .I(N__33569));
    LocalMux I__5921 (
            .O(N__33576),
            .I(N__33566));
    Sp12to4 I__5920 (
            .O(N__33569),
            .I(N__33563));
    Span4Mux_h I__5919 (
            .O(N__33566),
            .I(N__33560));
    Odrv12 I__5918 (
            .O(N__33563),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__5917 (
            .O(N__33560),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__5916 (
            .O(N__33555),
            .I(N__33552));
    LocalMux I__5915 (
            .O(N__33552),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    CascadeMux I__5914 (
            .O(N__33549),
            .I(N__33546));
    InMux I__5913 (
            .O(N__33546),
            .I(N__33541));
    InMux I__5912 (
            .O(N__33545),
            .I(N__33536));
    InMux I__5911 (
            .O(N__33544),
            .I(N__33536));
    LocalMux I__5910 (
            .O(N__33541),
            .I(N__33533));
    LocalMux I__5909 (
            .O(N__33536),
            .I(N__33530));
    Span4Mux_h I__5908 (
            .O(N__33533),
            .I(N__33526));
    Span4Mux_v I__5907 (
            .O(N__33530),
            .I(N__33523));
    InMux I__5906 (
            .O(N__33529),
            .I(N__33520));
    Odrv4 I__5905 (
            .O(N__33526),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__5904 (
            .O(N__33523),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__5903 (
            .O(N__33520),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    CascadeMux I__5902 (
            .O(N__33513),
            .I(N__33510));
    InMux I__5901 (
            .O(N__33510),
            .I(N__33505));
    InMux I__5900 (
            .O(N__33509),
            .I(N__33502));
    InMux I__5899 (
            .O(N__33508),
            .I(N__33499));
    LocalMux I__5898 (
            .O(N__33505),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__5897 (
            .O(N__33502),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__5896 (
            .O(N__33499),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__5895 (
            .O(N__33492),
            .I(N__33489));
    LocalMux I__5894 (
            .O(N__33489),
            .I(N__33486));
    Span4Mux_h I__5893 (
            .O(N__33486),
            .I(N__33483));
    Odrv4 I__5892 (
            .O(N__33483),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__5891 (
            .O(N__33480),
            .I(N__33477));
    LocalMux I__5890 (
            .O(N__33477),
            .I(N__33474));
    Span4Mux_v I__5889 (
            .O(N__33474),
            .I(N__33471));
    Odrv4 I__5888 (
            .O(N__33471),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ));
    ClkMux I__5887 (
            .O(N__33468),
            .I(N__33465));
    GlobalMux I__5886 (
            .O(N__33465),
            .I(N__33462));
    gio2CtrlBuf I__5885 (
            .O(N__33462),
            .I(delay_tr_input_c_g));
    InMux I__5884 (
            .O(N__33459),
            .I(N__33456));
    LocalMux I__5883 (
            .O(N__33456),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__5882 (
            .O(N__33453),
            .I(N__33449));
    CascadeMux I__5881 (
            .O(N__33452),
            .I(N__33446));
    InMux I__5880 (
            .O(N__33449),
            .I(N__33443));
    InMux I__5879 (
            .O(N__33446),
            .I(N__33440));
    LocalMux I__5878 (
            .O(N__33443),
            .I(N__33435));
    LocalMux I__5877 (
            .O(N__33440),
            .I(N__33432));
    InMux I__5876 (
            .O(N__33439),
            .I(N__33429));
    InMux I__5875 (
            .O(N__33438),
            .I(N__33426));
    Span12Mux_v I__5874 (
            .O(N__33435),
            .I(N__33423));
    Span12Mux_h I__5873 (
            .O(N__33432),
            .I(N__33416));
    LocalMux I__5872 (
            .O(N__33429),
            .I(N__33416));
    LocalMux I__5871 (
            .O(N__33426),
            .I(N__33416));
    Odrv12 I__5870 (
            .O(N__33423),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__5869 (
            .O(N__33416),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__5868 (
            .O(N__33411),
            .I(N__33406));
    InMux I__5867 (
            .O(N__33410),
            .I(N__33403));
    InMux I__5866 (
            .O(N__33409),
            .I(N__33400));
    LocalMux I__5865 (
            .O(N__33406),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__5864 (
            .O(N__33403),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__5863 (
            .O(N__33400),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__5862 (
            .O(N__33393),
            .I(N__33390));
    InMux I__5861 (
            .O(N__33390),
            .I(N__33387));
    LocalMux I__5860 (
            .O(N__33387),
            .I(N__33384));
    Span4Mux_v I__5859 (
            .O(N__33384),
            .I(N__33381));
    Odrv4 I__5858 (
            .O(N__33381),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__5857 (
            .O(N__33378),
            .I(N__33375));
    LocalMux I__5856 (
            .O(N__33375),
            .I(N__33371));
    InMux I__5855 (
            .O(N__33374),
            .I(N__33368));
    Span4Mux_h I__5854 (
            .O(N__33371),
            .I(N__33364));
    LocalMux I__5853 (
            .O(N__33368),
            .I(N__33361));
    InMux I__5852 (
            .O(N__33367),
            .I(N__33358));
    Span4Mux_v I__5851 (
            .O(N__33364),
            .I(N__33352));
    Span4Mux_h I__5850 (
            .O(N__33361),
            .I(N__33352));
    LocalMux I__5849 (
            .O(N__33358),
            .I(N__33349));
    InMux I__5848 (
            .O(N__33357),
            .I(N__33346));
    Span4Mux_v I__5847 (
            .O(N__33352),
            .I(N__33343));
    Span4Mux_v I__5846 (
            .O(N__33349),
            .I(N__33338));
    LocalMux I__5845 (
            .O(N__33346),
            .I(N__33338));
    Odrv4 I__5844 (
            .O(N__33343),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__5843 (
            .O(N__33338),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__5842 (
            .O(N__33333),
            .I(N__33329));
    CascadeMux I__5841 (
            .O(N__33332),
            .I(N__33325));
    LocalMux I__5840 (
            .O(N__33329),
            .I(N__33322));
    InMux I__5839 (
            .O(N__33328),
            .I(N__33319));
    InMux I__5838 (
            .O(N__33325),
            .I(N__33316));
    Span4Mux_v I__5837 (
            .O(N__33322),
            .I(N__33313));
    LocalMux I__5836 (
            .O(N__33319),
            .I(N__33310));
    LocalMux I__5835 (
            .O(N__33316),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__5834 (
            .O(N__33313),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__5833 (
            .O(N__33310),
            .I(\current_shift_inst.un4_control_input1_16 ));
    CascadeMux I__5832 (
            .O(N__33303),
            .I(N__33300));
    InMux I__5831 (
            .O(N__33300),
            .I(N__33297));
    LocalMux I__5830 (
            .O(N__33297),
            .I(N__33294));
    Span4Mux_v I__5829 (
            .O(N__33294),
            .I(N__33291));
    Span4Mux_h I__5828 (
            .O(N__33291),
            .I(N__33288));
    Odrv4 I__5827 (
            .O(N__33288),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__5826 (
            .O(N__33285),
            .I(N__33282));
    LocalMux I__5825 (
            .O(N__33282),
            .I(N__33277));
    CascadeMux I__5824 (
            .O(N__33281),
            .I(N__33274));
    InMux I__5823 (
            .O(N__33280),
            .I(N__33271));
    Span4Mux_h I__5822 (
            .O(N__33277),
            .I(N__33268));
    InMux I__5821 (
            .O(N__33274),
            .I(N__33265));
    LocalMux I__5820 (
            .O(N__33271),
            .I(N__33262));
    Odrv4 I__5819 (
            .O(N__33268),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__5818 (
            .O(N__33265),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__5817 (
            .O(N__33262),
            .I(\current_shift_inst.un4_control_input1_14 ));
    CascadeMux I__5816 (
            .O(N__33255),
            .I(N__33252));
    InMux I__5815 (
            .O(N__33252),
            .I(N__33249));
    LocalMux I__5814 (
            .O(N__33249),
            .I(N__33245));
    InMux I__5813 (
            .O(N__33248),
            .I(N__33242));
    Span4Mux_h I__5812 (
            .O(N__33245),
            .I(N__33238));
    LocalMux I__5811 (
            .O(N__33242),
            .I(N__33235));
    InMux I__5810 (
            .O(N__33241),
            .I(N__33232));
    Span4Mux_v I__5809 (
            .O(N__33238),
            .I(N__33226));
    Span4Mux_h I__5808 (
            .O(N__33235),
            .I(N__33226));
    LocalMux I__5807 (
            .O(N__33232),
            .I(N__33223));
    InMux I__5806 (
            .O(N__33231),
            .I(N__33220));
    Span4Mux_v I__5805 (
            .O(N__33226),
            .I(N__33217));
    Sp12to4 I__5804 (
            .O(N__33223),
            .I(N__33212));
    LocalMux I__5803 (
            .O(N__33220),
            .I(N__33212));
    Odrv4 I__5802 (
            .O(N__33217),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv12 I__5801 (
            .O(N__33212),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    CascadeMux I__5800 (
            .O(N__33207),
            .I(N__33204));
    InMux I__5799 (
            .O(N__33204),
            .I(N__33201));
    LocalMux I__5798 (
            .O(N__33201),
            .I(N__33198));
    Span4Mux_v I__5797 (
            .O(N__33198),
            .I(N__33195));
    Span4Mux_h I__5796 (
            .O(N__33195),
            .I(N__33192));
    Odrv4 I__5795 (
            .O(N__33192),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__5794 (
            .O(N__33189),
            .I(N__33186));
    LocalMux I__5793 (
            .O(N__33186),
            .I(N__33182));
    CascadeMux I__5792 (
            .O(N__33185),
            .I(N__33178));
    Span4Mux_h I__5791 (
            .O(N__33182),
            .I(N__33175));
    InMux I__5790 (
            .O(N__33181),
            .I(N__33172));
    InMux I__5789 (
            .O(N__33178),
            .I(N__33169));
    Odrv4 I__5788 (
            .O(N__33175),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__5787 (
            .O(N__33172),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__5786 (
            .O(N__33169),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__5785 (
            .O(N__33162),
            .I(N__33158));
    InMux I__5784 (
            .O(N__33161),
            .I(N__33155));
    LocalMux I__5783 (
            .O(N__33158),
            .I(N__33151));
    LocalMux I__5782 (
            .O(N__33155),
            .I(N__33148));
    InMux I__5781 (
            .O(N__33154),
            .I(N__33145));
    Span4Mux_v I__5780 (
            .O(N__33151),
            .I(N__33140));
    Span4Mux_v I__5779 (
            .O(N__33148),
            .I(N__33140));
    LocalMux I__5778 (
            .O(N__33145),
            .I(N__33137));
    Span4Mux_h I__5777 (
            .O(N__33140),
            .I(N__33133));
    Span4Mux_h I__5776 (
            .O(N__33137),
            .I(N__33130));
    InMux I__5775 (
            .O(N__33136),
            .I(N__33127));
    Odrv4 I__5774 (
            .O(N__33133),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    Odrv4 I__5773 (
            .O(N__33130),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__5772 (
            .O(N__33127),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__5771 (
            .O(N__33120),
            .I(N__33117));
    InMux I__5770 (
            .O(N__33117),
            .I(N__33114));
    LocalMux I__5769 (
            .O(N__33114),
            .I(N__33111));
    Span4Mux_v I__5768 (
            .O(N__33111),
            .I(N__33108));
    Odrv4 I__5767 (
            .O(N__33108),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt26 ));
    InMux I__5766 (
            .O(N__33105),
            .I(N__33101));
    CascadeMux I__5765 (
            .O(N__33104),
            .I(N__33097));
    LocalMux I__5764 (
            .O(N__33101),
            .I(N__33091));
    InMux I__5763 (
            .O(N__33100),
            .I(N__33086));
    InMux I__5762 (
            .O(N__33097),
            .I(N__33086));
    InMux I__5761 (
            .O(N__33096),
            .I(N__33083));
    InMux I__5760 (
            .O(N__33095),
            .I(N__33078));
    InMux I__5759 (
            .O(N__33094),
            .I(N__33078));
    Span4Mux_h I__5758 (
            .O(N__33091),
            .I(N__33075));
    LocalMux I__5757 (
            .O(N__33086),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__5756 (
            .O(N__33083),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__5755 (
            .O(N__33078),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__5754 (
            .O(N__33075),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__5753 (
            .O(N__33066),
            .I(N__33063));
    LocalMux I__5752 (
            .O(N__33063),
            .I(N__33060));
    Span4Mux_v I__5751 (
            .O(N__33060),
            .I(N__33057));
    Odrv4 I__5750 (
            .O(N__33057),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ));
    InMux I__5749 (
            .O(N__33054),
            .I(N__33051));
    LocalMux I__5748 (
            .O(N__33051),
            .I(N__33048));
    Span4Mux_v I__5747 (
            .O(N__33048),
            .I(N__33045));
    Odrv4 I__5746 (
            .O(N__33045),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ));
    InMux I__5745 (
            .O(N__33042),
            .I(N__33039));
    LocalMux I__5744 (
            .O(N__33039),
            .I(N__33036));
    Span4Mux_v I__5743 (
            .O(N__33036),
            .I(N__33033));
    Odrv4 I__5742 (
            .O(N__33033),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ));
    CascadeMux I__5741 (
            .O(N__33030),
            .I(N__33026));
    CascadeMux I__5740 (
            .O(N__33029),
            .I(N__33023));
    InMux I__5739 (
            .O(N__33026),
            .I(N__33018));
    InMux I__5738 (
            .O(N__33023),
            .I(N__33018));
    LocalMux I__5737 (
            .O(N__33018),
            .I(N__33015));
    Span4Mux_h I__5736 (
            .O(N__33015),
            .I(N__33012));
    Odrv4 I__5735 (
            .O(N__33012),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ));
    InMux I__5734 (
            .O(N__33009),
            .I(N__33006));
    LocalMux I__5733 (
            .O(N__33006),
            .I(N__33003));
    Span4Mux_v I__5732 (
            .O(N__33003),
            .I(N__33000));
    Span4Mux_h I__5731 (
            .O(N__33000),
            .I(N__32997));
    Span4Mux_h I__5730 (
            .O(N__32997),
            .I(N__32994));
    Odrv4 I__5729 (
            .O(N__32994),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ));
    InMux I__5728 (
            .O(N__32991),
            .I(N__32988));
    LocalMux I__5727 (
            .O(N__32988),
            .I(N__32985));
    Span4Mux_v I__5726 (
            .O(N__32985),
            .I(N__32982));
    Odrv4 I__5725 (
            .O(N__32982),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ));
    InMux I__5724 (
            .O(N__32979),
            .I(N__32976));
    LocalMux I__5723 (
            .O(N__32976),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt22 ));
    InMux I__5722 (
            .O(N__32973),
            .I(N__32968));
    InMux I__5721 (
            .O(N__32972),
            .I(N__32963));
    InMux I__5720 (
            .O(N__32971),
            .I(N__32963));
    LocalMux I__5719 (
            .O(N__32968),
            .I(N__32958));
    LocalMux I__5718 (
            .O(N__32963),
            .I(N__32958));
    Odrv4 I__5717 (
            .O(N__32958),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ));
    InMux I__5716 (
            .O(N__32955),
            .I(N__32950));
    InMux I__5715 (
            .O(N__32954),
            .I(N__32945));
    InMux I__5714 (
            .O(N__32953),
            .I(N__32945));
    LocalMux I__5713 (
            .O(N__32950),
            .I(N__32940));
    LocalMux I__5712 (
            .O(N__32945),
            .I(N__32940));
    Odrv4 I__5711 (
            .O(N__32940),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ));
    CascadeMux I__5710 (
            .O(N__32937),
            .I(N__32934));
    InMux I__5709 (
            .O(N__32934),
            .I(N__32931));
    LocalMux I__5708 (
            .O(N__32931),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ));
    InMux I__5707 (
            .O(N__32928),
            .I(N__32925));
    LocalMux I__5706 (
            .O(N__32925),
            .I(N__32922));
    Span4Mux_h I__5705 (
            .O(N__32922),
            .I(N__32919));
    Odrv4 I__5704 (
            .O(N__32919),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ));
    InMux I__5703 (
            .O(N__32916),
            .I(N__32913));
    LocalMux I__5702 (
            .O(N__32913),
            .I(N__32910));
    Odrv4 I__5701 (
            .O(N__32910),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ));
    InMux I__5700 (
            .O(N__32907),
            .I(N__32904));
    LocalMux I__5699 (
            .O(N__32904),
            .I(N__32901));
    Odrv4 I__5698 (
            .O(N__32901),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ));
    InMux I__5697 (
            .O(N__32898),
            .I(N__32892));
    InMux I__5696 (
            .O(N__32897),
            .I(N__32892));
    LocalMux I__5695 (
            .O(N__32892),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ));
    InMux I__5694 (
            .O(N__32889),
            .I(N__32883));
    InMux I__5693 (
            .O(N__32888),
            .I(N__32883));
    LocalMux I__5692 (
            .O(N__32883),
            .I(N__32880));
    Odrv4 I__5691 (
            .O(N__32880),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ));
    InMux I__5690 (
            .O(N__32877),
            .I(N__32873));
    InMux I__5689 (
            .O(N__32876),
            .I(N__32869));
    LocalMux I__5688 (
            .O(N__32873),
            .I(N__32866));
    InMux I__5687 (
            .O(N__32872),
            .I(N__32863));
    LocalMux I__5686 (
            .O(N__32869),
            .I(N__32860));
    Span4Mux_v I__5685 (
            .O(N__32866),
            .I(N__32857));
    LocalMux I__5684 (
            .O(N__32863),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    Odrv4 I__5683 (
            .O(N__32860),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    Odrv4 I__5682 (
            .O(N__32857),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    CascadeMux I__5681 (
            .O(N__32850),
            .I(N__32846));
    CascadeMux I__5680 (
            .O(N__32849),
            .I(N__32843));
    InMux I__5679 (
            .O(N__32846),
            .I(N__32839));
    InMux I__5678 (
            .O(N__32843),
            .I(N__32836));
    InMux I__5677 (
            .O(N__32842),
            .I(N__32833));
    LocalMux I__5676 (
            .O(N__32839),
            .I(N__32830));
    LocalMux I__5675 (
            .O(N__32836),
            .I(N__32827));
    LocalMux I__5674 (
            .O(N__32833),
            .I(N__32822));
    Span4Mux_v I__5673 (
            .O(N__32830),
            .I(N__32822));
    Odrv4 I__5672 (
            .O(N__32827),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ));
    Odrv4 I__5671 (
            .O(N__32822),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ));
    InMux I__5670 (
            .O(N__32817),
            .I(N__32810));
    InMux I__5669 (
            .O(N__32816),
            .I(N__32810));
    InMux I__5668 (
            .O(N__32815),
            .I(N__32807));
    LocalMux I__5667 (
            .O(N__32810),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__5666 (
            .O(N__32807),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__5665 (
            .O(N__32802),
            .I(N__32794));
    InMux I__5664 (
            .O(N__32801),
            .I(N__32789));
    InMux I__5663 (
            .O(N__32800),
            .I(N__32789));
    InMux I__5662 (
            .O(N__32799),
            .I(N__32784));
    InMux I__5661 (
            .O(N__32798),
            .I(N__32784));
    CascadeMux I__5660 (
            .O(N__32797),
            .I(N__32781));
    LocalMux I__5659 (
            .O(N__32794),
            .I(N__32778));
    LocalMux I__5658 (
            .O(N__32789),
            .I(N__32775));
    LocalMux I__5657 (
            .O(N__32784),
            .I(N__32772));
    InMux I__5656 (
            .O(N__32781),
            .I(N__32769));
    Span4Mux_v I__5655 (
            .O(N__32778),
            .I(N__32766));
    Span4Mux_v I__5654 (
            .O(N__32775),
            .I(N__32761));
    Span4Mux_v I__5653 (
            .O(N__32772),
            .I(N__32761));
    LocalMux I__5652 (
            .O(N__32769),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5651 (
            .O(N__32766),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5650 (
            .O(N__32761),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__5649 (
            .O(N__32754),
            .I(N__32751));
    LocalMux I__5648 (
            .O(N__32751),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ));
    InMux I__5647 (
            .O(N__32748),
            .I(N__32745));
    LocalMux I__5646 (
            .O(N__32745),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ));
    InMux I__5645 (
            .O(N__32742),
            .I(N__32739));
    LocalMux I__5644 (
            .O(N__32739),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ));
    InMux I__5643 (
            .O(N__32736),
            .I(N__32733));
    LocalMux I__5642 (
            .O(N__32733),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ));
    InMux I__5641 (
            .O(N__32730),
            .I(N__32727));
    LocalMux I__5640 (
            .O(N__32727),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ));
    CascadeMux I__5639 (
            .O(N__32724),
            .I(N__32721));
    InMux I__5638 (
            .O(N__32721),
            .I(N__32718));
    LocalMux I__5637 (
            .O(N__32718),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt20 ));
    InMux I__5636 (
            .O(N__32715),
            .I(N__32708));
    InMux I__5635 (
            .O(N__32714),
            .I(N__32708));
    InMux I__5634 (
            .O(N__32713),
            .I(N__32705));
    LocalMux I__5633 (
            .O(N__32708),
            .I(N__32702));
    LocalMux I__5632 (
            .O(N__32705),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ));
    Odrv4 I__5631 (
            .O(N__32702),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ));
    InMux I__5630 (
            .O(N__32697),
            .I(N__32690));
    InMux I__5629 (
            .O(N__32696),
            .I(N__32690));
    InMux I__5628 (
            .O(N__32695),
            .I(N__32687));
    LocalMux I__5627 (
            .O(N__32690),
            .I(N__32684));
    LocalMux I__5626 (
            .O(N__32687),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ));
    Odrv4 I__5625 (
            .O(N__32684),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ));
    InMux I__5624 (
            .O(N__32679),
            .I(N__32676));
    LocalMux I__5623 (
            .O(N__32676),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ));
    CascadeMux I__5622 (
            .O(N__32673),
            .I(N__32670));
    InMux I__5621 (
            .O(N__32670),
            .I(N__32667));
    LocalMux I__5620 (
            .O(N__32667),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ));
    InMux I__5619 (
            .O(N__32664),
            .I(N__32661));
    LocalMux I__5618 (
            .O(N__32661),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt20 ));
    InMux I__5617 (
            .O(N__32658),
            .I(N__32655));
    LocalMux I__5616 (
            .O(N__32655),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt22 ));
    CascadeMux I__5615 (
            .O(N__32652),
            .I(N__32649));
    InMux I__5614 (
            .O(N__32649),
            .I(N__32646));
    LocalMux I__5613 (
            .O(N__32646),
            .I(N__32643));
    Odrv4 I__5612 (
            .O(N__32643),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__5611 (
            .O(N__32640),
            .I(N__32637));
    InMux I__5610 (
            .O(N__32637),
            .I(N__32634));
    LocalMux I__5609 (
            .O(N__32634),
            .I(N__32631));
    Odrv4 I__5608 (
            .O(N__32631),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__5607 (
            .O(N__32628),
            .I(N__32625));
    LocalMux I__5606 (
            .O(N__32625),
            .I(N__32622));
    Odrv4 I__5605 (
            .O(N__32622),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt30 ));
    InMux I__5604 (
            .O(N__32619),
            .I(N__32616));
    LocalMux I__5603 (
            .O(N__32616),
            .I(N__32613));
    Odrv4 I__5602 (
            .O(N__32613),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt24 ));
    CEMux I__5601 (
            .O(N__32610),
            .I(N__32606));
    CEMux I__5600 (
            .O(N__32609),
            .I(N__32603));
    LocalMux I__5599 (
            .O(N__32606),
            .I(N__32599));
    LocalMux I__5598 (
            .O(N__32603),
            .I(N__32595));
    CEMux I__5597 (
            .O(N__32602),
            .I(N__32592));
    Span4Mux_h I__5596 (
            .O(N__32599),
            .I(N__32589));
    CEMux I__5595 (
            .O(N__32598),
            .I(N__32586));
    Span4Mux_h I__5594 (
            .O(N__32595),
            .I(N__32583));
    LocalMux I__5593 (
            .O(N__32592),
            .I(N__32580));
    Span4Mux_v I__5592 (
            .O(N__32589),
            .I(N__32577));
    LocalMux I__5591 (
            .O(N__32586),
            .I(N__32574));
    Span4Mux_v I__5590 (
            .O(N__32583),
            .I(N__32571));
    Span4Mux_h I__5589 (
            .O(N__32580),
            .I(N__32568));
    Span4Mux_v I__5588 (
            .O(N__32577),
            .I(N__32565));
    Span12Mux_v I__5587 (
            .O(N__32574),
            .I(N__32562));
    Sp12to4 I__5586 (
            .O(N__32571),
            .I(N__32557));
    Sp12to4 I__5585 (
            .O(N__32568),
            .I(N__32557));
    Odrv4 I__5584 (
            .O(N__32565),
            .I(\current_shift_inst.timer_s1.N_154_i ));
    Odrv12 I__5583 (
            .O(N__32562),
            .I(\current_shift_inst.timer_s1.N_154_i ));
    Odrv12 I__5582 (
            .O(N__32557),
            .I(\current_shift_inst.timer_s1.N_154_i ));
    CascadeMux I__5581 (
            .O(N__32550),
            .I(N__32547));
    InMux I__5580 (
            .O(N__32547),
            .I(N__32544));
    LocalMux I__5579 (
            .O(N__32544),
            .I(N__32541));
    Span4Mux_v I__5578 (
            .O(N__32541),
            .I(N__32538));
    Odrv4 I__5577 (
            .O(N__32538),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ));
    CascadeMux I__5576 (
            .O(N__32535),
            .I(N__32532));
    InMux I__5575 (
            .O(N__32532),
            .I(N__32529));
    LocalMux I__5574 (
            .O(N__32529),
            .I(N__32526));
    Odrv12 I__5573 (
            .O(N__32526),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt26 ));
    InMux I__5572 (
            .O(N__32523),
            .I(N__32520));
    LocalMux I__5571 (
            .O(N__32520),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__5570 (
            .O(N__32517),
            .I(bfn_11_28_0_));
    CascadeMux I__5569 (
            .O(N__32514),
            .I(N__32511));
    InMux I__5568 (
            .O(N__32511),
            .I(N__32508));
    LocalMux I__5567 (
            .O(N__32508),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt28 ));
    CascadeMux I__5566 (
            .O(N__32505),
            .I(N__32502));
    InMux I__5565 (
            .O(N__32502),
            .I(N__32499));
    LocalMux I__5564 (
            .O(N__32499),
            .I(\phase_controller_inst1.stoper_tr.counter_i_10 ));
    CascadeMux I__5563 (
            .O(N__32496),
            .I(N__32493));
    InMux I__5562 (
            .O(N__32493),
            .I(N__32490));
    LocalMux I__5561 (
            .O(N__32490),
            .I(N__32487));
    Odrv4 I__5560 (
            .O(N__32487),
            .I(\phase_controller_inst1.stoper_tr.counter_i_11 ));
    CascadeMux I__5559 (
            .O(N__32484),
            .I(N__32481));
    InMux I__5558 (
            .O(N__32481),
            .I(N__32478));
    LocalMux I__5557 (
            .O(N__32478),
            .I(N__32475));
    Odrv4 I__5556 (
            .O(N__32475),
            .I(\phase_controller_inst1.stoper_tr.counter_i_12 ));
    CascadeMux I__5555 (
            .O(N__32472),
            .I(N__32469));
    InMux I__5554 (
            .O(N__32469),
            .I(N__32466));
    LocalMux I__5553 (
            .O(N__32466),
            .I(N__32463));
    Odrv4 I__5552 (
            .O(N__32463),
            .I(\phase_controller_inst1.stoper_tr.counter_i_13 ));
    CascadeMux I__5551 (
            .O(N__32460),
            .I(N__32457));
    InMux I__5550 (
            .O(N__32457),
            .I(N__32454));
    LocalMux I__5549 (
            .O(N__32454),
            .I(N__32451));
    Odrv4 I__5548 (
            .O(N__32451),
            .I(\phase_controller_inst1.stoper_tr.counter_i_14 ));
    CascadeMux I__5547 (
            .O(N__32448),
            .I(N__32445));
    InMux I__5546 (
            .O(N__32445),
            .I(N__32442));
    LocalMux I__5545 (
            .O(N__32442),
            .I(\phase_controller_inst1.stoper_tr.counter_i_15 ));
    CascadeMux I__5544 (
            .O(N__32439),
            .I(N__32436));
    InMux I__5543 (
            .O(N__32436),
            .I(N__32433));
    LocalMux I__5542 (
            .O(N__32433),
            .I(\phase_controller_inst1.stoper_tr.counter_i_1 ));
    CascadeMux I__5541 (
            .O(N__32430),
            .I(N__32427));
    InMux I__5540 (
            .O(N__32427),
            .I(N__32424));
    LocalMux I__5539 (
            .O(N__32424),
            .I(\phase_controller_inst1.stoper_tr.counter_i_2 ));
    CascadeMux I__5538 (
            .O(N__32421),
            .I(N__32418));
    InMux I__5537 (
            .O(N__32418),
            .I(N__32415));
    LocalMux I__5536 (
            .O(N__32415),
            .I(\phase_controller_inst1.stoper_tr.counter_i_3 ));
    CascadeMux I__5535 (
            .O(N__32412),
            .I(N__32409));
    InMux I__5534 (
            .O(N__32409),
            .I(N__32406));
    LocalMux I__5533 (
            .O(N__32406),
            .I(N__32403));
    Odrv4 I__5532 (
            .O(N__32403),
            .I(\phase_controller_inst1.stoper_tr.counter_i_4 ));
    CascadeMux I__5531 (
            .O(N__32400),
            .I(N__32397));
    InMux I__5530 (
            .O(N__32397),
            .I(N__32394));
    LocalMux I__5529 (
            .O(N__32394),
            .I(\phase_controller_inst1.stoper_tr.counter_i_5 ));
    CascadeMux I__5528 (
            .O(N__32391),
            .I(N__32388));
    InMux I__5527 (
            .O(N__32388),
            .I(N__32385));
    LocalMux I__5526 (
            .O(N__32385),
            .I(N__32382));
    Odrv4 I__5525 (
            .O(N__32382),
            .I(\phase_controller_inst1.stoper_tr.counter_i_6 ));
    CascadeMux I__5524 (
            .O(N__32379),
            .I(N__32376));
    InMux I__5523 (
            .O(N__32376),
            .I(N__32373));
    LocalMux I__5522 (
            .O(N__32373),
            .I(\phase_controller_inst1.stoper_tr.counter_i_7 ));
    CascadeMux I__5521 (
            .O(N__32370),
            .I(N__32367));
    InMux I__5520 (
            .O(N__32367),
            .I(N__32364));
    LocalMux I__5519 (
            .O(N__32364),
            .I(\phase_controller_inst1.stoper_tr.counter_i_8 ));
    CascadeMux I__5518 (
            .O(N__32361),
            .I(N__32358));
    InMux I__5517 (
            .O(N__32358),
            .I(N__32355));
    LocalMux I__5516 (
            .O(N__32355),
            .I(\phase_controller_inst1.stoper_tr.counter_i_9 ));
    CascadeMux I__5515 (
            .O(N__32352),
            .I(N__32349));
    InMux I__5514 (
            .O(N__32349),
            .I(N__32346));
    LocalMux I__5513 (
            .O(N__32346),
            .I(N__32342));
    InMux I__5512 (
            .O(N__32345),
            .I(N__32339));
    Span4Mux_h I__5511 (
            .O(N__32342),
            .I(N__32335));
    LocalMux I__5510 (
            .O(N__32339),
            .I(N__32332));
    InMux I__5509 (
            .O(N__32338),
            .I(N__32329));
    Span4Mux_v I__5508 (
            .O(N__32335),
            .I(N__32323));
    Span4Mux_h I__5507 (
            .O(N__32332),
            .I(N__32323));
    LocalMux I__5506 (
            .O(N__32329),
            .I(N__32320));
    InMux I__5505 (
            .O(N__32328),
            .I(N__32317));
    Odrv4 I__5504 (
            .O(N__32323),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__5503 (
            .O(N__32320),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__5502 (
            .O(N__32317),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__5501 (
            .O(N__32310),
            .I(N__32307));
    LocalMux I__5500 (
            .O(N__32307),
            .I(N__32304));
    Odrv12 I__5499 (
            .O(N__32304),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__5498 (
            .O(N__32301),
            .I(N__32297));
    CascadeMux I__5497 (
            .O(N__32300),
            .I(N__32294));
    LocalMux I__5496 (
            .O(N__32297),
            .I(N__32290));
    InMux I__5495 (
            .O(N__32294),
            .I(N__32287));
    InMux I__5494 (
            .O(N__32293),
            .I(N__32284));
    Span4Mux_v I__5493 (
            .O(N__32290),
            .I(N__32277));
    LocalMux I__5492 (
            .O(N__32287),
            .I(N__32277));
    LocalMux I__5491 (
            .O(N__32284),
            .I(N__32277));
    Span4Mux_v I__5490 (
            .O(N__32277),
            .I(N__32273));
    InMux I__5489 (
            .O(N__32276),
            .I(N__32270));
    Odrv4 I__5488 (
            .O(N__32273),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__5487 (
            .O(N__32270),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__5486 (
            .O(N__32265),
            .I(N__32262));
    LocalMux I__5485 (
            .O(N__32262),
            .I(N__32259));
    Odrv12 I__5484 (
            .O(N__32259),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__5483 (
            .O(N__32256),
            .I(N__32253));
    LocalMux I__5482 (
            .O(N__32253),
            .I(N__32248));
    InMux I__5481 (
            .O(N__32252),
            .I(N__32245));
    InMux I__5480 (
            .O(N__32251),
            .I(N__32242));
    Span4Mux_v I__5479 (
            .O(N__32248),
            .I(N__32235));
    LocalMux I__5478 (
            .O(N__32245),
            .I(N__32235));
    LocalMux I__5477 (
            .O(N__32242),
            .I(N__32235));
    Span4Mux_v I__5476 (
            .O(N__32235),
            .I(N__32231));
    InMux I__5475 (
            .O(N__32234),
            .I(N__32228));
    Odrv4 I__5474 (
            .O(N__32231),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__5473 (
            .O(N__32228),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__5472 (
            .O(N__32223),
            .I(N__32220));
    LocalMux I__5471 (
            .O(N__32220),
            .I(N__32217));
    Span4Mux_v I__5470 (
            .O(N__32217),
            .I(N__32214));
    Odrv4 I__5469 (
            .O(N__32214),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    CascadeMux I__5468 (
            .O(N__32211),
            .I(N__32208));
    InMux I__5467 (
            .O(N__32208),
            .I(N__32205));
    LocalMux I__5466 (
            .O(N__32205),
            .I(N__32201));
    InMux I__5465 (
            .O(N__32204),
            .I(N__32198));
    Span4Mux_v I__5464 (
            .O(N__32201),
            .I(N__32192));
    LocalMux I__5463 (
            .O(N__32198),
            .I(N__32192));
    InMux I__5462 (
            .O(N__32197),
            .I(N__32189));
    Span4Mux_h I__5461 (
            .O(N__32192),
            .I(N__32186));
    LocalMux I__5460 (
            .O(N__32189),
            .I(N__32183));
    Span4Mux_v I__5459 (
            .O(N__32186),
            .I(N__32179));
    Span4Mux_v I__5458 (
            .O(N__32183),
            .I(N__32176));
    InMux I__5457 (
            .O(N__32182),
            .I(N__32173));
    Odrv4 I__5456 (
            .O(N__32179),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__5455 (
            .O(N__32176),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__5454 (
            .O(N__32173),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__5453 (
            .O(N__32166),
            .I(N__32163));
    LocalMux I__5452 (
            .O(N__32163),
            .I(N__32160));
    Odrv12 I__5451 (
            .O(N__32160),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    CascadeMux I__5450 (
            .O(N__32157),
            .I(N__32154));
    InMux I__5449 (
            .O(N__32154),
            .I(N__32151));
    LocalMux I__5448 (
            .O(N__32151),
            .I(N__32146));
    InMux I__5447 (
            .O(N__32150),
            .I(N__32141));
    InMux I__5446 (
            .O(N__32149),
            .I(N__32141));
    Span4Mux_v I__5445 (
            .O(N__32146),
            .I(N__32135));
    LocalMux I__5444 (
            .O(N__32141),
            .I(N__32135));
    InMux I__5443 (
            .O(N__32140),
            .I(N__32132));
    Span4Mux_v I__5442 (
            .O(N__32135),
            .I(N__32129));
    LocalMux I__5441 (
            .O(N__32132),
            .I(N__32126));
    Odrv4 I__5440 (
            .O(N__32129),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__5439 (
            .O(N__32126),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__5438 (
            .O(N__32121),
            .I(N__32118));
    LocalMux I__5437 (
            .O(N__32118),
            .I(N__32115));
    Span4Mux_v I__5436 (
            .O(N__32115),
            .I(N__32112));
    Span4Mux_v I__5435 (
            .O(N__32112),
            .I(N__32109));
    Odrv4 I__5434 (
            .O(N__32109),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__5433 (
            .O(N__32106),
            .I(N__32103));
    LocalMux I__5432 (
            .O(N__32103),
            .I(N__32099));
    InMux I__5431 (
            .O(N__32102),
            .I(N__32095));
    Span4Mux_h I__5430 (
            .O(N__32099),
            .I(N__32092));
    InMux I__5429 (
            .O(N__32098),
            .I(N__32089));
    LocalMux I__5428 (
            .O(N__32095),
            .I(N__32085));
    Span4Mux_v I__5427 (
            .O(N__32092),
            .I(N__32080));
    LocalMux I__5426 (
            .O(N__32089),
            .I(N__32080));
    InMux I__5425 (
            .O(N__32088),
            .I(N__32077));
    Span4Mux_v I__5424 (
            .O(N__32085),
            .I(N__32074));
    Span4Mux_v I__5423 (
            .O(N__32080),
            .I(N__32069));
    LocalMux I__5422 (
            .O(N__32077),
            .I(N__32069));
    Odrv4 I__5421 (
            .O(N__32074),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__5420 (
            .O(N__32069),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__5419 (
            .O(N__32064),
            .I(N__32061));
    LocalMux I__5418 (
            .O(N__32061),
            .I(N__32058));
    Sp12to4 I__5417 (
            .O(N__32058),
            .I(N__32055));
    Odrv12 I__5416 (
            .O(N__32055),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__5415 (
            .O(N__32052),
            .I(N__32049));
    LocalMux I__5414 (
            .O(N__32049),
            .I(\phase_controller_inst1.stoper_tr.counter_i_0 ));
    InMux I__5413 (
            .O(N__32046),
            .I(N__32043));
    LocalMux I__5412 (
            .O(N__32043),
            .I(N__32040));
    Span4Mux_h I__5411 (
            .O(N__32040),
            .I(N__32037));
    Span4Mux_h I__5410 (
            .O(N__32037),
            .I(N__32034));
    Span4Mux_v I__5409 (
            .O(N__32034),
            .I(N__32031));
    Odrv4 I__5408 (
            .O(N__32031),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    CascadeMux I__5407 (
            .O(N__32028),
            .I(N__32025));
    InMux I__5406 (
            .O(N__32025),
            .I(N__32022));
    LocalMux I__5405 (
            .O(N__32022),
            .I(N__32019));
    Span4Mux_h I__5404 (
            .O(N__32019),
            .I(N__32013));
    InMux I__5403 (
            .O(N__32018),
            .I(N__32008));
    InMux I__5402 (
            .O(N__32017),
            .I(N__32008));
    InMux I__5401 (
            .O(N__32016),
            .I(N__32005));
    Sp12to4 I__5400 (
            .O(N__32013),
            .I(N__32002));
    LocalMux I__5399 (
            .O(N__32008),
            .I(N__31999));
    LocalMux I__5398 (
            .O(N__32005),
            .I(N__31996));
    Span12Mux_v I__5397 (
            .O(N__32002),
            .I(N__31993));
    Span4Mux_h I__5396 (
            .O(N__31999),
            .I(N__31990));
    Odrv4 I__5395 (
            .O(N__31996),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv12 I__5394 (
            .O(N__31993),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__5393 (
            .O(N__31990),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__5392 (
            .O(N__31983),
            .I(bfn_11_22_0_));
    InMux I__5391 (
            .O(N__31980),
            .I(N__31977));
    LocalMux I__5390 (
            .O(N__31977),
            .I(N__31974));
    Span4Mux_h I__5389 (
            .O(N__31974),
            .I(N__31971));
    Span4Mux_h I__5388 (
            .O(N__31971),
            .I(N__31968));
    Odrv4 I__5387 (
            .O(N__31968),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    CascadeMux I__5386 (
            .O(N__31965),
            .I(N__31962));
    InMux I__5385 (
            .O(N__31962),
            .I(N__31959));
    LocalMux I__5384 (
            .O(N__31959),
            .I(N__31955));
    CascadeMux I__5383 (
            .O(N__31958),
            .I(N__31950));
    Span4Mux_v I__5382 (
            .O(N__31955),
            .I(N__31947));
    InMux I__5381 (
            .O(N__31954),
            .I(N__31944));
    InMux I__5380 (
            .O(N__31953),
            .I(N__31939));
    InMux I__5379 (
            .O(N__31950),
            .I(N__31939));
    Span4Mux_v I__5378 (
            .O(N__31947),
            .I(N__31936));
    LocalMux I__5377 (
            .O(N__31944),
            .I(N__31931));
    LocalMux I__5376 (
            .O(N__31939),
            .I(N__31931));
    Sp12to4 I__5375 (
            .O(N__31936),
            .I(N__31928));
    Span4Mux_h I__5374 (
            .O(N__31931),
            .I(N__31925));
    Odrv12 I__5373 (
            .O(N__31928),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__5372 (
            .O(N__31925),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__5371 (
            .O(N__31920),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__5370 (
            .O(N__31917),
            .I(N__31914));
    LocalMux I__5369 (
            .O(N__31914),
            .I(N__31911));
    Span4Mux_h I__5368 (
            .O(N__31911),
            .I(N__31908));
    Span4Mux_h I__5367 (
            .O(N__31908),
            .I(N__31905));
    Span4Mux_v I__5366 (
            .O(N__31905),
            .I(N__31902));
    Odrv4 I__5365 (
            .O(N__31902),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    CascadeMux I__5364 (
            .O(N__31899),
            .I(N__31896));
    InMux I__5363 (
            .O(N__31896),
            .I(N__31893));
    LocalMux I__5362 (
            .O(N__31893),
            .I(N__31890));
    Span4Mux_h I__5361 (
            .O(N__31890),
            .I(N__31887));
    Span4Mux_h I__5360 (
            .O(N__31887),
            .I(N__31883));
    InMux I__5359 (
            .O(N__31886),
            .I(N__31879));
    Sp12to4 I__5358 (
            .O(N__31883),
            .I(N__31875));
    InMux I__5357 (
            .O(N__31882),
            .I(N__31872));
    LocalMux I__5356 (
            .O(N__31879),
            .I(N__31869));
    InMux I__5355 (
            .O(N__31878),
            .I(N__31866));
    Span12Mux_v I__5354 (
            .O(N__31875),
            .I(N__31863));
    LocalMux I__5353 (
            .O(N__31872),
            .I(N__31858));
    Span4Mux_v I__5352 (
            .O(N__31869),
            .I(N__31858));
    LocalMux I__5351 (
            .O(N__31866),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__5350 (
            .O(N__31863),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__5349 (
            .O(N__31858),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__5348 (
            .O(N__31851),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__5347 (
            .O(N__31848),
            .I(N__31845));
    LocalMux I__5346 (
            .O(N__31845),
            .I(N__31842));
    Odrv12 I__5345 (
            .O(N__31842),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    CascadeMux I__5344 (
            .O(N__31839),
            .I(N__31836));
    InMux I__5343 (
            .O(N__31836),
            .I(N__31833));
    LocalMux I__5342 (
            .O(N__31833),
            .I(N__31830));
    Span4Mux_h I__5341 (
            .O(N__31830),
            .I(N__31827));
    Span4Mux_h I__5340 (
            .O(N__31827),
            .I(N__31821));
    CascadeMux I__5339 (
            .O(N__31826),
            .I(N__31818));
    InMux I__5338 (
            .O(N__31825),
            .I(N__31815));
    CascadeMux I__5337 (
            .O(N__31824),
            .I(N__31812));
    Span4Mux_v I__5336 (
            .O(N__31821),
            .I(N__31809));
    InMux I__5335 (
            .O(N__31818),
            .I(N__31806));
    LocalMux I__5334 (
            .O(N__31815),
            .I(N__31803));
    InMux I__5333 (
            .O(N__31812),
            .I(N__31800));
    Span4Mux_v I__5332 (
            .O(N__31809),
            .I(N__31795));
    LocalMux I__5331 (
            .O(N__31806),
            .I(N__31795));
    Span4Mux_v I__5330 (
            .O(N__31803),
            .I(N__31792));
    LocalMux I__5329 (
            .O(N__31800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__5328 (
            .O(N__31795),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__5327 (
            .O(N__31792),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__5326 (
            .O(N__31785),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__5325 (
            .O(N__31782),
            .I(N__31779));
    LocalMux I__5324 (
            .O(N__31779),
            .I(N__31776));
    Span4Mux_h I__5323 (
            .O(N__31776),
            .I(N__31773));
    Span4Mux_h I__5322 (
            .O(N__31773),
            .I(N__31770));
    Span4Mux_v I__5321 (
            .O(N__31770),
            .I(N__31767));
    Odrv4 I__5320 (
            .O(N__31767),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    CascadeMux I__5319 (
            .O(N__31764),
            .I(N__31761));
    InMux I__5318 (
            .O(N__31761),
            .I(N__31758));
    LocalMux I__5317 (
            .O(N__31758),
            .I(N__31753));
    InMux I__5316 (
            .O(N__31757),
            .I(N__31748));
    InMux I__5315 (
            .O(N__31756),
            .I(N__31748));
    Sp12to4 I__5314 (
            .O(N__31753),
            .I(N__31744));
    LocalMux I__5313 (
            .O(N__31748),
            .I(N__31741));
    InMux I__5312 (
            .O(N__31747),
            .I(N__31738));
    Span12Mux_v I__5311 (
            .O(N__31744),
            .I(N__31735));
    Span4Mux_h I__5310 (
            .O(N__31741),
            .I(N__31732));
    LocalMux I__5309 (
            .O(N__31738),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv12 I__5308 (
            .O(N__31735),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__5307 (
            .O(N__31732),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__5306 (
            .O(N__31725),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__5305 (
            .O(N__31722),
            .I(N__31719));
    LocalMux I__5304 (
            .O(N__31719),
            .I(N__31716));
    Odrv12 I__5303 (
            .O(N__31716),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    CascadeMux I__5302 (
            .O(N__31713),
            .I(N__31710));
    InMux I__5301 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__5300 (
            .O(N__31707),
            .I(N__31703));
    CascadeMux I__5299 (
            .O(N__31706),
            .I(N__31700));
    Span4Mux_h I__5298 (
            .O(N__31703),
            .I(N__31697));
    InMux I__5297 (
            .O(N__31700),
            .I(N__31694));
    Span4Mux_h I__5296 (
            .O(N__31697),
            .I(N__31691));
    LocalMux I__5295 (
            .O(N__31694),
            .I(N__31686));
    Span4Mux_v I__5294 (
            .O(N__31691),
            .I(N__31683));
    InMux I__5293 (
            .O(N__31690),
            .I(N__31680));
    InMux I__5292 (
            .O(N__31689),
            .I(N__31677));
    Span4Mux_h I__5291 (
            .O(N__31686),
            .I(N__31674));
    Span4Mux_v I__5290 (
            .O(N__31683),
            .I(N__31669));
    LocalMux I__5289 (
            .O(N__31680),
            .I(N__31669));
    LocalMux I__5288 (
            .O(N__31677),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5287 (
            .O(N__31674),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5286 (
            .O(N__31669),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__5285 (
            .O(N__31662),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__5284 (
            .O(N__31659),
            .I(N__31656));
    LocalMux I__5283 (
            .O(N__31656),
            .I(N__31644));
    InMux I__5282 (
            .O(N__31655),
            .I(N__31637));
    InMux I__5281 (
            .O(N__31654),
            .I(N__31626));
    InMux I__5280 (
            .O(N__31653),
            .I(N__31626));
    InMux I__5279 (
            .O(N__31652),
            .I(N__31626));
    InMux I__5278 (
            .O(N__31651),
            .I(N__31626));
    InMux I__5277 (
            .O(N__31650),
            .I(N__31617));
    InMux I__5276 (
            .O(N__31649),
            .I(N__31617));
    InMux I__5275 (
            .O(N__31648),
            .I(N__31617));
    InMux I__5274 (
            .O(N__31647),
            .I(N__31617));
    Span4Mux_v I__5273 (
            .O(N__31644),
            .I(N__31614));
    InMux I__5272 (
            .O(N__31643),
            .I(N__31610));
    InMux I__5271 (
            .O(N__31642),
            .I(N__31605));
    InMux I__5270 (
            .O(N__31641),
            .I(N__31605));
    InMux I__5269 (
            .O(N__31640),
            .I(N__31602));
    LocalMux I__5268 (
            .O(N__31637),
            .I(N__31599));
    InMux I__5267 (
            .O(N__31636),
            .I(N__31596));
    InMux I__5266 (
            .O(N__31635),
            .I(N__31579));
    LocalMux I__5265 (
            .O(N__31626),
            .I(N__31574));
    LocalMux I__5264 (
            .O(N__31617),
            .I(N__31574));
    Sp12to4 I__5263 (
            .O(N__31614),
            .I(N__31571));
    InMux I__5262 (
            .O(N__31613),
            .I(N__31568));
    LocalMux I__5261 (
            .O(N__31610),
            .I(N__31563));
    LocalMux I__5260 (
            .O(N__31605),
            .I(N__31563));
    LocalMux I__5259 (
            .O(N__31602),
            .I(N__31560));
    Span4Mux_v I__5258 (
            .O(N__31599),
            .I(N__31555));
    LocalMux I__5257 (
            .O(N__31596),
            .I(N__31555));
    InMux I__5256 (
            .O(N__31595),
            .I(N__31552));
    InMux I__5255 (
            .O(N__31594),
            .I(N__31545));
    InMux I__5254 (
            .O(N__31593),
            .I(N__31545));
    InMux I__5253 (
            .O(N__31592),
            .I(N__31545));
    InMux I__5252 (
            .O(N__31591),
            .I(N__31542));
    InMux I__5251 (
            .O(N__31590),
            .I(N__31535));
    InMux I__5250 (
            .O(N__31589),
            .I(N__31535));
    InMux I__5249 (
            .O(N__31588),
            .I(N__31535));
    InMux I__5248 (
            .O(N__31587),
            .I(N__31522));
    InMux I__5247 (
            .O(N__31586),
            .I(N__31522));
    InMux I__5246 (
            .O(N__31585),
            .I(N__31522));
    InMux I__5245 (
            .O(N__31584),
            .I(N__31522));
    InMux I__5244 (
            .O(N__31583),
            .I(N__31522));
    InMux I__5243 (
            .O(N__31582),
            .I(N__31522));
    LocalMux I__5242 (
            .O(N__31579),
            .I(N__31517));
    Span4Mux_v I__5241 (
            .O(N__31574),
            .I(N__31517));
    Span12Mux_h I__5240 (
            .O(N__31571),
            .I(N__31514));
    LocalMux I__5239 (
            .O(N__31568),
            .I(N__31505));
    Span4Mux_v I__5238 (
            .O(N__31563),
            .I(N__31505));
    Span4Mux_h I__5237 (
            .O(N__31560),
            .I(N__31505));
    Span4Mux_h I__5236 (
            .O(N__31555),
            .I(N__31505));
    LocalMux I__5235 (
            .O(N__31552),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__5234 (
            .O(N__31545),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__5233 (
            .O(N__31542),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__5232 (
            .O(N__31535),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__5231 (
            .O(N__31522),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__5230 (
            .O(N__31517),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__5229 (
            .O(N__31514),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__5228 (
            .O(N__31505),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__5227 (
            .O(N__31488),
            .I(N__31485));
    LocalMux I__5226 (
            .O(N__31485),
            .I(N__31482));
    Span4Mux_h I__5225 (
            .O(N__31482),
            .I(N__31479));
    Span4Mux_h I__5224 (
            .O(N__31479),
            .I(N__31476));
    Odrv4 I__5223 (
            .O(N__31476),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__5222 (
            .O(N__31473),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    IoInMux I__5221 (
            .O(N__31470),
            .I(N__31467));
    LocalMux I__5220 (
            .O(N__31467),
            .I(N__31464));
    Span4Mux_s3_v I__5219 (
            .O(N__31464),
            .I(N__31461));
    Span4Mux_h I__5218 (
            .O(N__31461),
            .I(N__31458));
    Span4Mux_v I__5217 (
            .O(N__31458),
            .I(N__31455));
    Odrv4 I__5216 (
            .O(N__31455),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__5215 (
            .O(N__31452),
            .I(N__31449));
    LocalMux I__5214 (
            .O(N__31449),
            .I(N__31446));
    Odrv12 I__5213 (
            .O(N__31446),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__5212 (
            .O(N__31443),
            .I(N__31440));
    InMux I__5211 (
            .O(N__31440),
            .I(N__31437));
    LocalMux I__5210 (
            .O(N__31437),
            .I(N__31433));
    CascadeMux I__5209 (
            .O(N__31436),
            .I(N__31430));
    Span4Mux_v I__5208 (
            .O(N__31433),
            .I(N__31426));
    InMux I__5207 (
            .O(N__31430),
            .I(N__31423));
    InMux I__5206 (
            .O(N__31429),
            .I(N__31420));
    Sp12to4 I__5205 (
            .O(N__31426),
            .I(N__31416));
    LocalMux I__5204 (
            .O(N__31423),
            .I(N__31413));
    LocalMux I__5203 (
            .O(N__31420),
            .I(N__31410));
    InMux I__5202 (
            .O(N__31419),
            .I(N__31407));
    Span12Mux_h I__5201 (
            .O(N__31416),
            .I(N__31404));
    Span4Mux_h I__5200 (
            .O(N__31413),
            .I(N__31399));
    Span4Mux_h I__5199 (
            .O(N__31410),
            .I(N__31399));
    LocalMux I__5198 (
            .O(N__31407),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv12 I__5197 (
            .O(N__31404),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__5196 (
            .O(N__31399),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__5195 (
            .O(N__31392),
            .I(bfn_11_21_0_));
    InMux I__5194 (
            .O(N__31389),
            .I(N__31386));
    LocalMux I__5193 (
            .O(N__31386),
            .I(N__31383));
    Span4Mux_h I__5192 (
            .O(N__31383),
            .I(N__31380));
    Span4Mux_h I__5191 (
            .O(N__31380),
            .I(N__31377));
    Odrv4 I__5190 (
            .O(N__31377),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    CascadeMux I__5189 (
            .O(N__31374),
            .I(N__31371));
    InMux I__5188 (
            .O(N__31371),
            .I(N__31368));
    LocalMux I__5187 (
            .O(N__31368),
            .I(N__31365));
    Span4Mux_h I__5186 (
            .O(N__31365),
            .I(N__31362));
    Span4Mux_h I__5185 (
            .O(N__31362),
            .I(N__31357));
    InMux I__5184 (
            .O(N__31361),
            .I(N__31354));
    InMux I__5183 (
            .O(N__31360),
            .I(N__31351));
    Span4Mux_v I__5182 (
            .O(N__31357),
            .I(N__31345));
    LocalMux I__5181 (
            .O(N__31354),
            .I(N__31345));
    LocalMux I__5180 (
            .O(N__31351),
            .I(N__31342));
    InMux I__5179 (
            .O(N__31350),
            .I(N__31339));
    Span4Mux_v I__5178 (
            .O(N__31345),
            .I(N__31336));
    Odrv4 I__5177 (
            .O(N__31342),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__5176 (
            .O(N__31339),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__5175 (
            .O(N__31336),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__5174 (
            .O(N__31329),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__5173 (
            .O(N__31326),
            .I(N__31323));
    LocalMux I__5172 (
            .O(N__31323),
            .I(N__31320));
    Span4Mux_h I__5171 (
            .O(N__31320),
            .I(N__31317));
    Span4Mux_h I__5170 (
            .O(N__31317),
            .I(N__31314));
    Span4Mux_v I__5169 (
            .O(N__31314),
            .I(N__31311));
    Odrv4 I__5168 (
            .O(N__31311),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    CascadeMux I__5167 (
            .O(N__31308),
            .I(N__31304));
    CascadeMux I__5166 (
            .O(N__31307),
            .I(N__31300));
    InMux I__5165 (
            .O(N__31304),
            .I(N__31297));
    InMux I__5164 (
            .O(N__31303),
            .I(N__31293));
    InMux I__5163 (
            .O(N__31300),
            .I(N__31290));
    LocalMux I__5162 (
            .O(N__31297),
            .I(N__31287));
    InMux I__5161 (
            .O(N__31296),
            .I(N__31284));
    LocalMux I__5160 (
            .O(N__31293),
            .I(N__31281));
    LocalMux I__5159 (
            .O(N__31290),
            .I(N__31278));
    Span12Mux_h I__5158 (
            .O(N__31287),
            .I(N__31275));
    LocalMux I__5157 (
            .O(N__31284),
            .I(N__31272));
    Span4Mux_v I__5156 (
            .O(N__31281),
            .I(N__31267));
    Span4Mux_v I__5155 (
            .O(N__31278),
            .I(N__31267));
    Odrv12 I__5154 (
            .O(N__31275),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__5153 (
            .O(N__31272),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__5152 (
            .O(N__31267),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__5151 (
            .O(N__31260),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__5150 (
            .O(N__31257),
            .I(N__31254));
    LocalMux I__5149 (
            .O(N__31254),
            .I(N__31251));
    Span4Mux_h I__5148 (
            .O(N__31251),
            .I(N__31248));
    Span4Mux_h I__5147 (
            .O(N__31248),
            .I(N__31245));
    Odrv4 I__5146 (
            .O(N__31245),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__5145 (
            .O(N__31242),
            .I(N__31239));
    InMux I__5144 (
            .O(N__31239),
            .I(N__31236));
    LocalMux I__5143 (
            .O(N__31236),
            .I(N__31233));
    Span4Mux_v I__5142 (
            .O(N__31233),
            .I(N__31230));
    Span4Mux_h I__5141 (
            .O(N__31230),
            .I(N__31224));
    CascadeMux I__5140 (
            .O(N__31229),
            .I(N__31221));
    InMux I__5139 (
            .O(N__31228),
            .I(N__31218));
    InMux I__5138 (
            .O(N__31227),
            .I(N__31215));
    Span4Mux_h I__5137 (
            .O(N__31224),
            .I(N__31212));
    InMux I__5136 (
            .O(N__31221),
            .I(N__31209));
    LocalMux I__5135 (
            .O(N__31218),
            .I(N__31206));
    LocalMux I__5134 (
            .O(N__31215),
            .I(N__31203));
    Span4Mux_v I__5133 (
            .O(N__31212),
            .I(N__31200));
    LocalMux I__5132 (
            .O(N__31209),
            .I(N__31193));
    Span4Mux_h I__5131 (
            .O(N__31206),
            .I(N__31193));
    Span4Mux_h I__5130 (
            .O(N__31203),
            .I(N__31193));
    Odrv4 I__5129 (
            .O(N__31200),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__5128 (
            .O(N__31193),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__5127 (
            .O(N__31188),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__5126 (
            .O(N__31185),
            .I(N__31182));
    LocalMux I__5125 (
            .O(N__31182),
            .I(N__31179));
    Span4Mux_v I__5124 (
            .O(N__31179),
            .I(N__31176));
    Odrv4 I__5123 (
            .O(N__31176),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__5122 (
            .O(N__31173),
            .I(N__31170));
    InMux I__5121 (
            .O(N__31170),
            .I(N__31167));
    LocalMux I__5120 (
            .O(N__31167),
            .I(N__31164));
    Span4Mux_h I__5119 (
            .O(N__31164),
            .I(N__31161));
    Span4Mux_h I__5118 (
            .O(N__31161),
            .I(N__31158));
    Span4Mux_v I__5117 (
            .O(N__31158),
            .I(N__31152));
    InMux I__5116 (
            .O(N__31157),
            .I(N__31147));
    InMux I__5115 (
            .O(N__31156),
            .I(N__31147));
    InMux I__5114 (
            .O(N__31155),
            .I(N__31144));
    Span4Mux_v I__5113 (
            .O(N__31152),
            .I(N__31139));
    LocalMux I__5112 (
            .O(N__31147),
            .I(N__31139));
    LocalMux I__5111 (
            .O(N__31144),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__5110 (
            .O(N__31139),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__5109 (
            .O(N__31134),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__5108 (
            .O(N__31131),
            .I(N__31128));
    LocalMux I__5107 (
            .O(N__31128),
            .I(N__31125));
    Span12Mux_h I__5106 (
            .O(N__31125),
            .I(N__31122));
    Odrv12 I__5105 (
            .O(N__31122),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__5104 (
            .O(N__31119),
            .I(N__31116));
    InMux I__5103 (
            .O(N__31116),
            .I(N__31111));
    InMux I__5102 (
            .O(N__31115),
            .I(N__31108));
    InMux I__5101 (
            .O(N__31114),
            .I(N__31105));
    LocalMux I__5100 (
            .O(N__31111),
            .I(N__31102));
    LocalMux I__5099 (
            .O(N__31108),
            .I(N__31098));
    LocalMux I__5098 (
            .O(N__31105),
            .I(N__31095));
    Span12Mux_v I__5097 (
            .O(N__31102),
            .I(N__31092));
    InMux I__5096 (
            .O(N__31101),
            .I(N__31089));
    Span4Mux_h I__5095 (
            .O(N__31098),
            .I(N__31084));
    Span4Mux_h I__5094 (
            .O(N__31095),
            .I(N__31084));
    Odrv12 I__5093 (
            .O(N__31092),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__5092 (
            .O(N__31089),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5091 (
            .O(N__31084),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__5090 (
            .O(N__31077),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__5089 (
            .O(N__31074),
            .I(N__31071));
    LocalMux I__5088 (
            .O(N__31071),
            .I(N__31068));
    Span4Mux_h I__5087 (
            .O(N__31068),
            .I(N__31065));
    Odrv4 I__5086 (
            .O(N__31065),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__5085 (
            .O(N__31062),
            .I(N__31059));
    InMux I__5084 (
            .O(N__31059),
            .I(N__31056));
    LocalMux I__5083 (
            .O(N__31056),
            .I(N__31053));
    Span4Mux_v I__5082 (
            .O(N__31053),
            .I(N__31050));
    Span4Mux_v I__5081 (
            .O(N__31050),
            .I(N__31046));
    CascadeMux I__5080 (
            .O(N__31049),
            .I(N__31043));
    Span4Mux_v I__5079 (
            .O(N__31046),
            .I(N__31038));
    InMux I__5078 (
            .O(N__31043),
            .I(N__31033));
    InMux I__5077 (
            .O(N__31042),
            .I(N__31033));
    InMux I__5076 (
            .O(N__31041),
            .I(N__31030));
    Span4Mux_h I__5075 (
            .O(N__31038),
            .I(N__31025));
    LocalMux I__5074 (
            .O(N__31033),
            .I(N__31025));
    LocalMux I__5073 (
            .O(N__31030),
            .I(N__31020));
    Span4Mux_h I__5072 (
            .O(N__31025),
            .I(N__31020));
    Odrv4 I__5071 (
            .O(N__31020),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__5070 (
            .O(N__31017),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__5069 (
            .O(N__31014),
            .I(N__31011));
    LocalMux I__5068 (
            .O(N__31011),
            .I(N__31008));
    Span4Mux_h I__5067 (
            .O(N__31008),
            .I(N__31005));
    Span4Mux_h I__5066 (
            .O(N__31005),
            .I(N__31002));
    Odrv4 I__5065 (
            .O(N__31002),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__5064 (
            .O(N__30999),
            .I(N__30996));
    InMux I__5063 (
            .O(N__30996),
            .I(N__30993));
    LocalMux I__5062 (
            .O(N__30993),
            .I(N__30990));
    Span4Mux_v I__5061 (
            .O(N__30990),
            .I(N__30986));
    CascadeMux I__5060 (
            .O(N__30989),
            .I(N__30983));
    Sp12to4 I__5059 (
            .O(N__30986),
            .I(N__30978));
    InMux I__5058 (
            .O(N__30983),
            .I(N__30973));
    InMux I__5057 (
            .O(N__30982),
            .I(N__30973));
    InMux I__5056 (
            .O(N__30981),
            .I(N__30970));
    Span12Mux_h I__5055 (
            .O(N__30978),
            .I(N__30967));
    LocalMux I__5054 (
            .O(N__30973),
            .I(N__30964));
    LocalMux I__5053 (
            .O(N__30970),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__5052 (
            .O(N__30967),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__5051 (
            .O(N__30964),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__5050 (
            .O(N__30957),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__5049 (
            .O(N__30954),
            .I(N__30951));
    LocalMux I__5048 (
            .O(N__30951),
            .I(N__30948));
    Span4Mux_h I__5047 (
            .O(N__30948),
            .I(N__30945));
    Odrv4 I__5046 (
            .O(N__30945),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__5045 (
            .O(N__30942),
            .I(N__30939));
    InMux I__5044 (
            .O(N__30939),
            .I(N__30936));
    LocalMux I__5043 (
            .O(N__30936),
            .I(N__30933));
    Span4Mux_h I__5042 (
            .O(N__30933),
            .I(N__30930));
    Span4Mux_h I__5041 (
            .O(N__30930),
            .I(N__30924));
    InMux I__5040 (
            .O(N__30929),
            .I(N__30921));
    CascadeMux I__5039 (
            .O(N__30928),
            .I(N__30918));
    InMux I__5038 (
            .O(N__30927),
            .I(N__30915));
    Sp12to4 I__5037 (
            .O(N__30924),
            .I(N__30910));
    LocalMux I__5036 (
            .O(N__30921),
            .I(N__30910));
    InMux I__5035 (
            .O(N__30918),
            .I(N__30907));
    LocalMux I__5034 (
            .O(N__30915),
            .I(N__30904));
    Span12Mux_v I__5033 (
            .O(N__30910),
            .I(N__30901));
    LocalMux I__5032 (
            .O(N__30907),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__5031 (
            .O(N__30904),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__5030 (
            .O(N__30901),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__5029 (
            .O(N__30894),
            .I(bfn_11_20_0_));
    InMux I__5028 (
            .O(N__30891),
            .I(N__30888));
    LocalMux I__5027 (
            .O(N__30888),
            .I(N__30885));
    Span4Mux_h I__5026 (
            .O(N__30885),
            .I(N__30882));
    Span4Mux_h I__5025 (
            .O(N__30882),
            .I(N__30879));
    Span4Mux_v I__5024 (
            .O(N__30879),
            .I(N__30876));
    Odrv4 I__5023 (
            .O(N__30876),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__5022 (
            .O(N__30873),
            .I(N__30870));
    InMux I__5021 (
            .O(N__30870),
            .I(N__30867));
    LocalMux I__5020 (
            .O(N__30867),
            .I(N__30864));
    Span4Mux_v I__5019 (
            .O(N__30864),
            .I(N__30861));
    Span4Mux_h I__5018 (
            .O(N__30861),
            .I(N__30857));
    CascadeMux I__5017 (
            .O(N__30860),
            .I(N__30854));
    Span4Mux_h I__5016 (
            .O(N__30857),
            .I(N__30849));
    InMux I__5015 (
            .O(N__30854),
            .I(N__30846));
    InMux I__5014 (
            .O(N__30853),
            .I(N__30843));
    InMux I__5013 (
            .O(N__30852),
            .I(N__30840));
    Span4Mux_v I__5012 (
            .O(N__30849),
            .I(N__30835));
    LocalMux I__5011 (
            .O(N__30846),
            .I(N__30835));
    LocalMux I__5010 (
            .O(N__30843),
            .I(N__30830));
    LocalMux I__5009 (
            .O(N__30840),
            .I(N__30830));
    Odrv4 I__5008 (
            .O(N__30835),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__5007 (
            .O(N__30830),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__5006 (
            .O(N__30825),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__5005 (
            .O(N__30822),
            .I(N__30819));
    LocalMux I__5004 (
            .O(N__30819),
            .I(N__30816));
    Span4Mux_v I__5003 (
            .O(N__30816),
            .I(N__30813));
    Span4Mux_v I__5002 (
            .O(N__30813),
            .I(N__30810));
    Odrv4 I__5001 (
            .O(N__30810),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__5000 (
            .O(N__30807),
            .I(N__30804));
    InMux I__4999 (
            .O(N__30804),
            .I(N__30801));
    LocalMux I__4998 (
            .O(N__30801),
            .I(N__30798));
    Span4Mux_h I__4997 (
            .O(N__30798),
            .I(N__30795));
    Span4Mux_h I__4996 (
            .O(N__30795),
            .I(N__30790));
    CascadeMux I__4995 (
            .O(N__30794),
            .I(N__30787));
    InMux I__4994 (
            .O(N__30793),
            .I(N__30784));
    Span4Mux_v I__4993 (
            .O(N__30790),
            .I(N__30781));
    InMux I__4992 (
            .O(N__30787),
            .I(N__30778));
    LocalMux I__4991 (
            .O(N__30784),
            .I(N__30775));
    Span4Mux_v I__4990 (
            .O(N__30781),
            .I(N__30771));
    LocalMux I__4989 (
            .O(N__30778),
            .I(N__30766));
    Span4Mux_h I__4988 (
            .O(N__30775),
            .I(N__30766));
    InMux I__4987 (
            .O(N__30774),
            .I(N__30763));
    Odrv4 I__4986 (
            .O(N__30771),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__4985 (
            .O(N__30766),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__4984 (
            .O(N__30763),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__4983 (
            .O(N__30756),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__4982 (
            .O(N__30753),
            .I(N__30750));
    LocalMux I__4981 (
            .O(N__30750),
            .I(N__30747));
    Span4Mux_v I__4980 (
            .O(N__30747),
            .I(N__30744));
    Span4Mux_h I__4979 (
            .O(N__30744),
            .I(N__30741));
    Odrv4 I__4978 (
            .O(N__30741),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__4977 (
            .O(N__30738),
            .I(N__30735));
    InMux I__4976 (
            .O(N__30735),
            .I(N__30732));
    LocalMux I__4975 (
            .O(N__30732),
            .I(N__30728));
    CascadeMux I__4974 (
            .O(N__30731),
            .I(N__30724));
    Span4Mux_v I__4973 (
            .O(N__30728),
            .I(N__30720));
    InMux I__4972 (
            .O(N__30727),
            .I(N__30717));
    InMux I__4971 (
            .O(N__30724),
            .I(N__30714));
    InMux I__4970 (
            .O(N__30723),
            .I(N__30711));
    Span4Mux_h I__4969 (
            .O(N__30720),
            .I(N__30708));
    LocalMux I__4968 (
            .O(N__30717),
            .I(N__30705));
    LocalMux I__4967 (
            .O(N__30714),
            .I(N__30702));
    LocalMux I__4966 (
            .O(N__30711),
            .I(N__30699));
    Span4Mux_h I__4965 (
            .O(N__30708),
            .I(N__30694));
    Span4Mux_h I__4964 (
            .O(N__30705),
            .I(N__30694));
    Odrv12 I__4963 (
            .O(N__30702),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__4962 (
            .O(N__30699),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__4961 (
            .O(N__30694),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__4960 (
            .O(N__30687),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__4959 (
            .O(N__30684),
            .I(N__30681));
    LocalMux I__4958 (
            .O(N__30681),
            .I(N__30678));
    Span4Mux_v I__4957 (
            .O(N__30678),
            .I(N__30675));
    Span4Mux_v I__4956 (
            .O(N__30675),
            .I(N__30672));
    Odrv4 I__4955 (
            .O(N__30672),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__4954 (
            .O(N__30669),
            .I(N__30666));
    InMux I__4953 (
            .O(N__30666),
            .I(N__30663));
    LocalMux I__4952 (
            .O(N__30663),
            .I(N__30660));
    Span4Mux_v I__4951 (
            .O(N__30660),
            .I(N__30657));
    Sp12to4 I__4950 (
            .O(N__30657),
            .I(N__30652));
    InMux I__4949 (
            .O(N__30656),
            .I(N__30648));
    InMux I__4948 (
            .O(N__30655),
            .I(N__30645));
    Span12Mux_h I__4947 (
            .O(N__30652),
            .I(N__30642));
    InMux I__4946 (
            .O(N__30651),
            .I(N__30639));
    LocalMux I__4945 (
            .O(N__30648),
            .I(N__30636));
    LocalMux I__4944 (
            .O(N__30645),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv12 I__4943 (
            .O(N__30642),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__4942 (
            .O(N__30639),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__4941 (
            .O(N__30636),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__4940 (
            .O(N__30627),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__4939 (
            .O(N__30624),
            .I(N__30621));
    LocalMux I__4938 (
            .O(N__30621),
            .I(N__30618));
    Span4Mux_v I__4937 (
            .O(N__30618),
            .I(N__30615));
    Span4Mux_h I__4936 (
            .O(N__30615),
            .I(N__30612));
    Odrv4 I__4935 (
            .O(N__30612),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__4934 (
            .O(N__30609),
            .I(N__30606));
    InMux I__4933 (
            .O(N__30606),
            .I(N__30603));
    LocalMux I__4932 (
            .O(N__30603),
            .I(N__30599));
    InMux I__4931 (
            .O(N__30602),
            .I(N__30594));
    Span12Mux_v I__4930 (
            .O(N__30599),
            .I(N__30591));
    InMux I__4929 (
            .O(N__30598),
            .I(N__30588));
    InMux I__4928 (
            .O(N__30597),
            .I(N__30585));
    LocalMux I__4927 (
            .O(N__30594),
            .I(N__30582));
    Odrv12 I__4926 (
            .O(N__30591),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__4925 (
            .O(N__30588),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__4924 (
            .O(N__30585),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4923 (
            .O(N__30582),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__4922 (
            .O(N__30573),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__4921 (
            .O(N__30570),
            .I(N__30567));
    LocalMux I__4920 (
            .O(N__30567),
            .I(N__30564));
    Span4Mux_v I__4919 (
            .O(N__30564),
            .I(N__30561));
    Span4Mux_v I__4918 (
            .O(N__30561),
            .I(N__30558));
    Odrv4 I__4917 (
            .O(N__30558),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__4916 (
            .O(N__30555),
            .I(N__30552));
    InMux I__4915 (
            .O(N__30552),
            .I(N__30549));
    LocalMux I__4914 (
            .O(N__30549),
            .I(N__30544));
    CascadeMux I__4913 (
            .O(N__30548),
            .I(N__30541));
    InMux I__4912 (
            .O(N__30547),
            .I(N__30537));
    Span4Mux_v I__4911 (
            .O(N__30544),
            .I(N__30534));
    InMux I__4910 (
            .O(N__30541),
            .I(N__30531));
    InMux I__4909 (
            .O(N__30540),
            .I(N__30528));
    LocalMux I__4908 (
            .O(N__30537),
            .I(N__30525));
    Span4Mux_h I__4907 (
            .O(N__30534),
            .I(N__30522));
    LocalMux I__4906 (
            .O(N__30531),
            .I(N__30519));
    LocalMux I__4905 (
            .O(N__30528),
            .I(N__30516));
    Span4Mux_v I__4904 (
            .O(N__30525),
            .I(N__30513));
    Span4Mux_h I__4903 (
            .O(N__30522),
            .I(N__30508));
    Span4Mux_v I__4902 (
            .O(N__30519),
            .I(N__30508));
    Span4Mux_v I__4901 (
            .O(N__30516),
            .I(N__30505));
    Odrv4 I__4900 (
            .O(N__30513),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4899 (
            .O(N__30508),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4898 (
            .O(N__30505),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__4897 (
            .O(N__30498),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__4896 (
            .O(N__30495),
            .I(N__30492));
    LocalMux I__4895 (
            .O(N__30492),
            .I(N__30489));
    Span12Mux_v I__4894 (
            .O(N__30489),
            .I(N__30486));
    Odrv12 I__4893 (
            .O(N__30486),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    CascadeMux I__4892 (
            .O(N__30483),
            .I(N__30479));
    CascadeMux I__4891 (
            .O(N__30482),
            .I(N__30475));
    InMux I__4890 (
            .O(N__30479),
            .I(N__30472));
    InMux I__4889 (
            .O(N__30478),
            .I(N__30469));
    InMux I__4888 (
            .O(N__30475),
            .I(N__30466));
    LocalMux I__4887 (
            .O(N__30472),
            .I(N__30463));
    LocalMux I__4886 (
            .O(N__30469),
            .I(N__30459));
    LocalMux I__4885 (
            .O(N__30466),
            .I(N__30456));
    Span12Mux_v I__4884 (
            .O(N__30463),
            .I(N__30453));
    InMux I__4883 (
            .O(N__30462),
            .I(N__30450));
    Span4Mux_v I__4882 (
            .O(N__30459),
            .I(N__30445));
    Span4Mux_h I__4881 (
            .O(N__30456),
            .I(N__30445));
    Odrv12 I__4880 (
            .O(N__30453),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__4879 (
            .O(N__30450),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__4878 (
            .O(N__30445),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__4877 (
            .O(N__30438),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__4876 (
            .O(N__30435),
            .I(N__30432));
    LocalMux I__4875 (
            .O(N__30432),
            .I(N__30428));
    InMux I__4874 (
            .O(N__30431),
            .I(N__30424));
    Span12Mux_h I__4873 (
            .O(N__30428),
            .I(N__30421));
    InMux I__4872 (
            .O(N__30427),
            .I(N__30418));
    LocalMux I__4871 (
            .O(N__30424),
            .I(N__30415));
    Odrv12 I__4870 (
            .O(N__30421),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__4869 (
            .O(N__30418),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__4868 (
            .O(N__30415),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    CascadeMux I__4867 (
            .O(N__30408),
            .I(N__30405));
    InMux I__4866 (
            .O(N__30405),
            .I(N__30402));
    LocalMux I__4865 (
            .O(N__30402),
            .I(N__30399));
    Span4Mux_h I__4864 (
            .O(N__30399),
            .I(N__30396));
    Odrv4 I__4863 (
            .O(N__30396),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__4862 (
            .O(N__30393),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__4861 (
            .O(N__30390),
            .I(N__30387));
    LocalMux I__4860 (
            .O(N__30387),
            .I(N__30384));
    Span4Mux_h I__4859 (
            .O(N__30384),
            .I(N__30381));
    Span4Mux_h I__4858 (
            .O(N__30381),
            .I(N__30378));
    Odrv4 I__4857 (
            .O(N__30378),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__4856 (
            .O(N__30375),
            .I(N__30372));
    InMux I__4855 (
            .O(N__30372),
            .I(N__30369));
    LocalMux I__4854 (
            .O(N__30369),
            .I(N__30365));
    CascadeMux I__4853 (
            .O(N__30368),
            .I(N__30362));
    Span4Mux_v I__4852 (
            .O(N__30365),
            .I(N__30359));
    InMux I__4851 (
            .O(N__30362),
            .I(N__30356));
    Span4Mux_h I__4850 (
            .O(N__30359),
            .I(N__30353));
    LocalMux I__4849 (
            .O(N__30356),
            .I(N__30348));
    Span4Mux_h I__4848 (
            .O(N__30353),
            .I(N__30345));
    InMux I__4847 (
            .O(N__30352),
            .I(N__30342));
    InMux I__4846 (
            .O(N__30351),
            .I(N__30339));
    Span4Mux_h I__4845 (
            .O(N__30348),
            .I(N__30334));
    Span4Mux_v I__4844 (
            .O(N__30345),
            .I(N__30334));
    LocalMux I__4843 (
            .O(N__30342),
            .I(N__30331));
    LocalMux I__4842 (
            .O(N__30339),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__4841 (
            .O(N__30334),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__4840 (
            .O(N__30331),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__4839 (
            .O(N__30324),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__4838 (
            .O(N__30321),
            .I(N__30318));
    LocalMux I__4837 (
            .O(N__30318),
            .I(N__30315));
    Span4Mux_v I__4836 (
            .O(N__30315),
            .I(N__30312));
    Odrv4 I__4835 (
            .O(N__30312),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__4834 (
            .O(N__30309),
            .I(N__30306));
    InMux I__4833 (
            .O(N__30306),
            .I(N__30303));
    LocalMux I__4832 (
            .O(N__30303),
            .I(N__30300));
    Span4Mux_v I__4831 (
            .O(N__30300),
            .I(N__30297));
    Sp12to4 I__4830 (
            .O(N__30297),
            .I(N__30291));
    InMux I__4829 (
            .O(N__30296),
            .I(N__30288));
    InMux I__4828 (
            .O(N__30295),
            .I(N__30285));
    InMux I__4827 (
            .O(N__30294),
            .I(N__30282));
    Span12Mux_h I__4826 (
            .O(N__30291),
            .I(N__30279));
    LocalMux I__4825 (
            .O(N__30288),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__4824 (
            .O(N__30285),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__4823 (
            .O(N__30282),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__4822 (
            .O(N__30279),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__4821 (
            .O(N__30270),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__4820 (
            .O(N__30267),
            .I(N__30264));
    LocalMux I__4819 (
            .O(N__30264),
            .I(N__30261));
    Span4Mux_v I__4818 (
            .O(N__30261),
            .I(N__30258));
    Span4Mux_v I__4817 (
            .O(N__30258),
            .I(N__30255));
    Odrv4 I__4816 (
            .O(N__30255),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__4815 (
            .O(N__30252),
            .I(N__30249));
    InMux I__4814 (
            .O(N__30249),
            .I(N__30246));
    LocalMux I__4813 (
            .O(N__30246),
            .I(N__30243));
    Span4Mux_h I__4812 (
            .O(N__30243),
            .I(N__30240));
    Span4Mux_h I__4811 (
            .O(N__30240),
            .I(N__30236));
    InMux I__4810 (
            .O(N__30239),
            .I(N__30233));
    Span4Mux_h I__4809 (
            .O(N__30236),
            .I(N__30229));
    LocalMux I__4808 (
            .O(N__30233),
            .I(N__30225));
    InMux I__4807 (
            .O(N__30232),
            .I(N__30222));
    Sp12to4 I__4806 (
            .O(N__30229),
            .I(N__30219));
    InMux I__4805 (
            .O(N__30228),
            .I(N__30216));
    Span4Mux_h I__4804 (
            .O(N__30225),
            .I(N__30213));
    LocalMux I__4803 (
            .O(N__30222),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv12 I__4802 (
            .O(N__30219),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__4801 (
            .O(N__30216),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__4800 (
            .O(N__30213),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__4799 (
            .O(N__30204),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__4798 (
            .O(N__30201),
            .I(N__30198));
    LocalMux I__4797 (
            .O(N__30198),
            .I(N__30195));
    Span4Mux_v I__4796 (
            .O(N__30195),
            .I(N__30192));
    Span4Mux_v I__4795 (
            .O(N__30192),
            .I(N__30189));
    Odrv4 I__4794 (
            .O(N__30189),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__4793 (
            .O(N__30186),
            .I(N__30183));
    InMux I__4792 (
            .O(N__30183),
            .I(N__30180));
    LocalMux I__4791 (
            .O(N__30180),
            .I(N__30177));
    Span4Mux_v I__4790 (
            .O(N__30177),
            .I(N__30174));
    Sp12to4 I__4789 (
            .O(N__30174),
            .I(N__30168));
    InMux I__4788 (
            .O(N__30173),
            .I(N__30165));
    InMux I__4787 (
            .O(N__30172),
            .I(N__30162));
    InMux I__4786 (
            .O(N__30171),
            .I(N__30159));
    Span12Mux_h I__4785 (
            .O(N__30168),
            .I(N__30156));
    LocalMux I__4784 (
            .O(N__30165),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4783 (
            .O(N__30162),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4782 (
            .O(N__30159),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv12 I__4781 (
            .O(N__30156),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__4780 (
            .O(N__30147),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__4779 (
            .O(N__30144),
            .I(N__30141));
    LocalMux I__4778 (
            .O(N__30141),
            .I(N__30138));
    Span4Mux_v I__4777 (
            .O(N__30138),
            .I(N__30135));
    Span4Mux_h I__4776 (
            .O(N__30135),
            .I(N__30132));
    Odrv4 I__4775 (
            .O(N__30132),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__4774 (
            .O(N__30129),
            .I(N__30126));
    InMux I__4773 (
            .O(N__30126),
            .I(N__30123));
    LocalMux I__4772 (
            .O(N__30123),
            .I(N__30120));
    Span4Mux_v I__4771 (
            .O(N__30120),
            .I(N__30117));
    Span4Mux_h I__4770 (
            .O(N__30117),
            .I(N__30114));
    Span4Mux_h I__4769 (
            .O(N__30114),
            .I(N__30110));
    InMux I__4768 (
            .O(N__30113),
            .I(N__30107));
    Span4Mux_v I__4767 (
            .O(N__30110),
            .I(N__30100));
    LocalMux I__4766 (
            .O(N__30107),
            .I(N__30100));
    InMux I__4765 (
            .O(N__30106),
            .I(N__30097));
    InMux I__4764 (
            .O(N__30105),
            .I(N__30094));
    Span4Mux_v I__4763 (
            .O(N__30100),
            .I(N__30091));
    LocalMux I__4762 (
            .O(N__30097),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__4761 (
            .O(N__30094),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__4760 (
            .O(N__30091),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__4759 (
            .O(N__30084),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__4758 (
            .O(N__30081),
            .I(N__30078));
    LocalMux I__4757 (
            .O(N__30078),
            .I(N__30075));
    Odrv12 I__4756 (
            .O(N__30075),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__4755 (
            .O(N__30072),
            .I(N__30069));
    InMux I__4754 (
            .O(N__30069),
            .I(N__30066));
    LocalMux I__4753 (
            .O(N__30066),
            .I(N__30063));
    Span4Mux_v I__4752 (
            .O(N__30063),
            .I(N__30060));
    Sp12to4 I__4751 (
            .O(N__30060),
            .I(N__30054));
    InMux I__4750 (
            .O(N__30059),
            .I(N__30051));
    InMux I__4749 (
            .O(N__30058),
            .I(N__30048));
    InMux I__4748 (
            .O(N__30057),
            .I(N__30045));
    Span12Mux_v I__4747 (
            .O(N__30054),
            .I(N__30042));
    LocalMux I__4746 (
            .O(N__30051),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__4745 (
            .O(N__30048),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__4744 (
            .O(N__30045),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv12 I__4743 (
            .O(N__30042),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__4742 (
            .O(N__30033),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    CascadeMux I__4741 (
            .O(N__30030),
            .I(N__30027));
    InMux I__4740 (
            .O(N__30027),
            .I(N__30024));
    LocalMux I__4739 (
            .O(N__30024),
            .I(N__30019));
    InMux I__4738 (
            .O(N__30023),
            .I(N__30016));
    InMux I__4737 (
            .O(N__30022),
            .I(N__30013));
    Span4Mux_v I__4736 (
            .O(N__30019),
            .I(N__30008));
    LocalMux I__4735 (
            .O(N__30016),
            .I(N__30008));
    LocalMux I__4734 (
            .O(N__30013),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__4733 (
            .O(N__30008),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__4732 (
            .O(N__30003),
            .I(bfn_11_18_0_));
    InMux I__4731 (
            .O(N__30000),
            .I(N__29997));
    LocalMux I__4730 (
            .O(N__29997),
            .I(N__29994));
    Span4Mux_h I__4729 (
            .O(N__29994),
            .I(N__29991));
    Span4Mux_v I__4728 (
            .O(N__29991),
            .I(N__29988));
    Odrv4 I__4727 (
            .O(N__29988),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__4726 (
            .O(N__29985),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__4725 (
            .O(N__29982),
            .I(N__29979));
    LocalMux I__4724 (
            .O(N__29979),
            .I(N__29975));
    CascadeMux I__4723 (
            .O(N__29978),
            .I(N__29972));
    Span4Mux_h I__4722 (
            .O(N__29975),
            .I(N__29968));
    InMux I__4721 (
            .O(N__29972),
            .I(N__29965));
    InMux I__4720 (
            .O(N__29971),
            .I(N__29962));
    Odrv4 I__4719 (
            .O(N__29968),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__4718 (
            .O(N__29965),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__4717 (
            .O(N__29962),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__4716 (
            .O(N__29955),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__4715 (
            .O(N__29952),
            .I(N__29949));
    LocalMux I__4714 (
            .O(N__29949),
            .I(N__29946));
    Span4Mux_h I__4713 (
            .O(N__29946),
            .I(N__29941));
    InMux I__4712 (
            .O(N__29945),
            .I(N__29938));
    InMux I__4711 (
            .O(N__29944),
            .I(N__29935));
    Span4Mux_v I__4710 (
            .O(N__29941),
            .I(N__29930));
    LocalMux I__4709 (
            .O(N__29938),
            .I(N__29930));
    LocalMux I__4708 (
            .O(N__29935),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__4707 (
            .O(N__29930),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__4706 (
            .O(N__29925),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__4705 (
            .O(N__29922),
            .I(N__29918));
    InMux I__4704 (
            .O(N__29921),
            .I(N__29914));
    LocalMux I__4703 (
            .O(N__29918),
            .I(N__29911));
    InMux I__4702 (
            .O(N__29917),
            .I(N__29908));
    LocalMux I__4701 (
            .O(N__29914),
            .I(N__29905));
    Span4Mux_v I__4700 (
            .O(N__29911),
            .I(N__29900));
    LocalMux I__4699 (
            .O(N__29908),
            .I(N__29900));
    Odrv12 I__4698 (
            .O(N__29905),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__4697 (
            .O(N__29900),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__4696 (
            .O(N__29895),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__4695 (
            .O(N__29892),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__4694 (
            .O(N__29889),
            .I(N__29885));
    InMux I__4693 (
            .O(N__29888),
            .I(N__29882));
    InMux I__4692 (
            .O(N__29885),
            .I(N__29876));
    LocalMux I__4691 (
            .O(N__29882),
            .I(N__29873));
    CascadeMux I__4690 (
            .O(N__29881),
            .I(N__29870));
    InMux I__4689 (
            .O(N__29880),
            .I(N__29865));
    InMux I__4688 (
            .O(N__29879),
            .I(N__29865));
    LocalMux I__4687 (
            .O(N__29876),
            .I(N__29860));
    Span4Mux_v I__4686 (
            .O(N__29873),
            .I(N__29860));
    InMux I__4685 (
            .O(N__29870),
            .I(N__29857));
    LocalMux I__4684 (
            .O(N__29865),
            .I(N__29854));
    Sp12to4 I__4683 (
            .O(N__29860),
            .I(N__29849));
    LocalMux I__4682 (
            .O(N__29857),
            .I(N__29849));
    Span12Mux_v I__4681 (
            .O(N__29854),
            .I(N__29844));
    Span12Mux_h I__4680 (
            .O(N__29849),
            .I(N__29844));
    Odrv12 I__4679 (
            .O(N__29844),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__4678 (
            .O(N__29841),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__4677 (
            .O(N__29838),
            .I(N__29835));
    LocalMux I__4676 (
            .O(N__29835),
            .I(N__29832));
    Span4Mux_v I__4675 (
            .O(N__29832),
            .I(N__29829));
    Odrv4 I__4674 (
            .O(N__29829),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__4673 (
            .O(N__29826),
            .I(N__29823));
    LocalMux I__4672 (
            .O(N__29823),
            .I(N__29819));
    InMux I__4671 (
            .O(N__29822),
            .I(N__29815));
    Span4Mux_h I__4670 (
            .O(N__29819),
            .I(N__29812));
    InMux I__4669 (
            .O(N__29818),
            .I(N__29809));
    LocalMux I__4668 (
            .O(N__29815),
            .I(N__29806));
    Odrv4 I__4667 (
            .O(N__29812),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__4666 (
            .O(N__29809),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__4665 (
            .O(N__29806),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__4664 (
            .O(N__29799),
            .I(N__29796));
    InMux I__4663 (
            .O(N__29796),
            .I(N__29793));
    LocalMux I__4662 (
            .O(N__29793),
            .I(N__29790));
    Span4Mux_h I__4661 (
            .O(N__29790),
            .I(N__29787));
    Odrv4 I__4660 (
            .O(N__29787),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__4659 (
            .O(N__29784),
            .I(N__29781));
    LocalMux I__4658 (
            .O(N__29781),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__4657 (
            .O(N__29778),
            .I(N__29775));
    LocalMux I__4656 (
            .O(N__29775),
            .I(N__29771));
    InMux I__4655 (
            .O(N__29774),
            .I(N__29767));
    Span4Mux_h I__4654 (
            .O(N__29771),
            .I(N__29764));
    InMux I__4653 (
            .O(N__29770),
            .I(N__29761));
    LocalMux I__4652 (
            .O(N__29767),
            .I(N__29758));
    Odrv4 I__4651 (
            .O(N__29764),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__4650 (
            .O(N__29761),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__4649 (
            .O(N__29758),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__4648 (
            .O(N__29751),
            .I(bfn_11_17_0_));
    InMux I__4647 (
            .O(N__29748),
            .I(N__29745));
    LocalMux I__4646 (
            .O(N__29745),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__4645 (
            .O(N__29742),
            .I(N__29739));
    LocalMux I__4644 (
            .O(N__29739),
            .I(N__29735));
    InMux I__4643 (
            .O(N__29738),
            .I(N__29732));
    Span4Mux_v I__4642 (
            .O(N__29735),
            .I(N__29728));
    LocalMux I__4641 (
            .O(N__29732),
            .I(N__29725));
    InMux I__4640 (
            .O(N__29731),
            .I(N__29722));
    Span4Mux_h I__4639 (
            .O(N__29728),
            .I(N__29717));
    Span4Mux_h I__4638 (
            .O(N__29725),
            .I(N__29717));
    LocalMux I__4637 (
            .O(N__29722),
            .I(N__29714));
    Odrv4 I__4636 (
            .O(N__29717),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__4635 (
            .O(N__29714),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__4634 (
            .O(N__29709),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__4633 (
            .O(N__29706),
            .I(N__29703));
    LocalMux I__4632 (
            .O(N__29703),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__4631 (
            .O(N__29700),
            .I(N__29696));
    InMux I__4630 (
            .O(N__29699),
            .I(N__29693));
    LocalMux I__4629 (
            .O(N__29696),
            .I(N__29690));
    LocalMux I__4628 (
            .O(N__29693),
            .I(N__29686));
    Span4Mux_h I__4627 (
            .O(N__29690),
            .I(N__29683));
    InMux I__4626 (
            .O(N__29689),
            .I(N__29680));
    Span4Mux_h I__4625 (
            .O(N__29686),
            .I(N__29677));
    Span4Mux_v I__4624 (
            .O(N__29683),
            .I(N__29672));
    LocalMux I__4623 (
            .O(N__29680),
            .I(N__29672));
    Odrv4 I__4622 (
            .O(N__29677),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__4621 (
            .O(N__29672),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__4620 (
            .O(N__29667),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__4619 (
            .O(N__29664),
            .I(N__29661));
    LocalMux I__4618 (
            .O(N__29661),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__4617 (
            .O(N__29658),
            .I(N__29654));
    CascadeMux I__4616 (
            .O(N__29657),
            .I(N__29651));
    LocalMux I__4615 (
            .O(N__29654),
            .I(N__29647));
    InMux I__4614 (
            .O(N__29651),
            .I(N__29644));
    InMux I__4613 (
            .O(N__29650),
            .I(N__29641));
    Span4Mux_h I__4612 (
            .O(N__29647),
            .I(N__29636));
    LocalMux I__4611 (
            .O(N__29644),
            .I(N__29636));
    LocalMux I__4610 (
            .O(N__29641),
            .I(N__29633));
    Odrv4 I__4609 (
            .O(N__29636),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__4608 (
            .O(N__29633),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__4607 (
            .O(N__29628),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__4606 (
            .O(N__29625),
            .I(N__29622));
    LocalMux I__4605 (
            .O(N__29622),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    CascadeMux I__4604 (
            .O(N__29619),
            .I(N__29615));
    InMux I__4603 (
            .O(N__29618),
            .I(N__29612));
    InMux I__4602 (
            .O(N__29615),
            .I(N__29608));
    LocalMux I__4601 (
            .O(N__29612),
            .I(N__29605));
    InMux I__4600 (
            .O(N__29611),
            .I(N__29602));
    LocalMux I__4599 (
            .O(N__29608),
            .I(N__29599));
    Span4Mux_v I__4598 (
            .O(N__29605),
            .I(N__29594));
    LocalMux I__4597 (
            .O(N__29602),
            .I(N__29594));
    Odrv4 I__4596 (
            .O(N__29599),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__4595 (
            .O(N__29594),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__4594 (
            .O(N__29589),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__4593 (
            .O(N__29586),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__4592 (
            .O(N__29583),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    CascadeMux I__4591 (
            .O(N__29580),
            .I(N__29577));
    InMux I__4590 (
            .O(N__29577),
            .I(N__29573));
    InMux I__4589 (
            .O(N__29576),
            .I(N__29570));
    LocalMux I__4588 (
            .O(N__29573),
            .I(N__29567));
    LocalMux I__4587 (
            .O(N__29570),
            .I(N__29563));
    Span4Mux_v I__4586 (
            .O(N__29567),
            .I(N__29560));
    InMux I__4585 (
            .O(N__29566),
            .I(N__29557));
    Odrv12 I__4584 (
            .O(N__29563),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__4583 (
            .O(N__29560),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__4582 (
            .O(N__29557),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__4581 (
            .O(N__29550),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    CascadeMux I__4580 (
            .O(N__29547),
            .I(N__29544));
    InMux I__4579 (
            .O(N__29544),
            .I(N__29541));
    LocalMux I__4578 (
            .O(N__29541),
            .I(N__29538));
    Odrv4 I__4577 (
            .O(N__29538),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__4576 (
            .O(N__29535),
            .I(N__29531));
    InMux I__4575 (
            .O(N__29534),
            .I(N__29528));
    LocalMux I__4574 (
            .O(N__29531),
            .I(N__29524));
    LocalMux I__4573 (
            .O(N__29528),
            .I(N__29521));
    InMux I__4572 (
            .O(N__29527),
            .I(N__29518));
    Span4Mux_v I__4571 (
            .O(N__29524),
            .I(N__29511));
    Span4Mux_v I__4570 (
            .O(N__29521),
            .I(N__29511));
    LocalMux I__4569 (
            .O(N__29518),
            .I(N__29511));
    Odrv4 I__4568 (
            .O(N__29511),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__4567 (
            .O(N__29508),
            .I(bfn_11_16_0_));
    InMux I__4566 (
            .O(N__29505),
            .I(N__29502));
    LocalMux I__4565 (
            .O(N__29502),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__4564 (
            .O(N__29499),
            .I(N__29495));
    InMux I__4563 (
            .O(N__29498),
            .I(N__29492));
    LocalMux I__4562 (
            .O(N__29495),
            .I(N__29489));
    LocalMux I__4561 (
            .O(N__29492),
            .I(N__29486));
    Span4Mux_v I__4560 (
            .O(N__29489),
            .I(N__29483));
    Span4Mux_h I__4559 (
            .O(N__29486),
            .I(N__29479));
    Span4Mux_h I__4558 (
            .O(N__29483),
            .I(N__29476));
    InMux I__4557 (
            .O(N__29482),
            .I(N__29473));
    Odrv4 I__4556 (
            .O(N__29479),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__4555 (
            .O(N__29476),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__4554 (
            .O(N__29473),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__4553 (
            .O(N__29466),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__4552 (
            .O(N__29463),
            .I(N__29460));
    LocalMux I__4551 (
            .O(N__29460),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__4550 (
            .O(N__29457),
            .I(N__29453));
    InMux I__4549 (
            .O(N__29456),
            .I(N__29450));
    LocalMux I__4548 (
            .O(N__29453),
            .I(N__29447));
    LocalMux I__4547 (
            .O(N__29450),
            .I(N__29443));
    Span4Mux_v I__4546 (
            .O(N__29447),
            .I(N__29440));
    InMux I__4545 (
            .O(N__29446),
            .I(N__29437));
    Span4Mux_h I__4544 (
            .O(N__29443),
            .I(N__29434));
    Span4Mux_v I__4543 (
            .O(N__29440),
            .I(N__29429));
    LocalMux I__4542 (
            .O(N__29437),
            .I(N__29429));
    Odrv4 I__4541 (
            .O(N__29434),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__4540 (
            .O(N__29429),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__4539 (
            .O(N__29424),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__4538 (
            .O(N__29421),
            .I(N__29418));
    LocalMux I__4537 (
            .O(N__29418),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__4536 (
            .O(N__29415),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__4535 (
            .O(N__29412),
            .I(N__29409));
    LocalMux I__4534 (
            .O(N__29409),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__4533 (
            .O(N__29406),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__4532 (
            .O(N__29403),
            .I(N__29400));
    LocalMux I__4531 (
            .O(N__29400),
            .I(N__29397));
    Odrv4 I__4530 (
            .O(N__29397),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__4529 (
            .O(N__29394),
            .I(N__29391));
    LocalMux I__4528 (
            .O(N__29391),
            .I(N__29386));
    InMux I__4527 (
            .O(N__29390),
            .I(N__29381));
    InMux I__4526 (
            .O(N__29389),
            .I(N__29381));
    Odrv4 I__4525 (
            .O(N__29386),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__4524 (
            .O(N__29381),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__4523 (
            .O(N__29376),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__4522 (
            .O(N__29373),
            .I(N__29370));
    LocalMux I__4521 (
            .O(N__29370),
            .I(N__29367));
    Odrv4 I__4520 (
            .O(N__29367),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__4519 (
            .O(N__29364),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__4518 (
            .O(N__29361),
            .I(N__29358));
    LocalMux I__4517 (
            .O(N__29358),
            .I(N__29353));
    InMux I__4516 (
            .O(N__29357),
            .I(N__29348));
    InMux I__4515 (
            .O(N__29356),
            .I(N__29348));
    Span4Mux_v I__4514 (
            .O(N__29353),
            .I(N__29345));
    LocalMux I__4513 (
            .O(N__29348),
            .I(N__29342));
    Odrv4 I__4512 (
            .O(N__29345),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv12 I__4511 (
            .O(N__29342),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__4510 (
            .O(N__29337),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    CascadeMux I__4509 (
            .O(N__29334),
            .I(N__29331));
    InMux I__4508 (
            .O(N__29331),
            .I(N__29326));
    InMux I__4507 (
            .O(N__29330),
            .I(N__29323));
    InMux I__4506 (
            .O(N__29329),
            .I(N__29320));
    LocalMux I__4505 (
            .O(N__29326),
            .I(N__29317));
    LocalMux I__4504 (
            .O(N__29323),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__4503 (
            .O(N__29320),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__4502 (
            .O(N__29317),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__4501 (
            .O(N__29310),
            .I(N__29306));
    InMux I__4500 (
            .O(N__29309),
            .I(N__29303));
    InMux I__4499 (
            .O(N__29306),
            .I(N__29300));
    LocalMux I__4498 (
            .O(N__29303),
            .I(N__29296));
    LocalMux I__4497 (
            .O(N__29300),
            .I(N__29293));
    InMux I__4496 (
            .O(N__29299),
            .I(N__29290));
    Span4Mux_v I__4495 (
            .O(N__29296),
            .I(N__29283));
    Span4Mux_v I__4494 (
            .O(N__29293),
            .I(N__29283));
    LocalMux I__4493 (
            .O(N__29290),
            .I(N__29283));
    Odrv4 I__4492 (
            .O(N__29283),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__4491 (
            .O(N__29280),
            .I(N__29277));
    LocalMux I__4490 (
            .O(N__29277),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__4489 (
            .O(N__29274),
            .I(N__29271));
    LocalMux I__4488 (
            .O(N__29271),
            .I(N__29267));
    InMux I__4487 (
            .O(N__29270),
            .I(N__29264));
    Span4Mux_v I__4486 (
            .O(N__29267),
            .I(N__29260));
    LocalMux I__4485 (
            .O(N__29264),
            .I(N__29257));
    InMux I__4484 (
            .O(N__29263),
            .I(N__29254));
    Odrv4 I__4483 (
            .O(N__29260),
            .I(\current_shift_inst.un4_control_input1_3 ));
    Odrv4 I__4482 (
            .O(N__29257),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__4481 (
            .O(N__29254),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__4480 (
            .O(N__29247),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__4479 (
            .O(N__29244),
            .I(N__29241));
    LocalMux I__4478 (
            .O(N__29241),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    CascadeMux I__4477 (
            .O(N__29238),
            .I(N__29235));
    InMux I__4476 (
            .O(N__29235),
            .I(N__29232));
    LocalMux I__4475 (
            .O(N__29232),
            .I(N__29228));
    InMux I__4474 (
            .O(N__29231),
            .I(N__29225));
    Span4Mux_h I__4473 (
            .O(N__29228),
            .I(N__29221));
    LocalMux I__4472 (
            .O(N__29225),
            .I(N__29218));
    InMux I__4471 (
            .O(N__29224),
            .I(N__29215));
    Odrv4 I__4470 (
            .O(N__29221),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__4469 (
            .O(N__29218),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__4468 (
            .O(N__29215),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__4467 (
            .O(N__29208),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__4466 (
            .O(N__29205),
            .I(N__29202));
    LocalMux I__4465 (
            .O(N__29202),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    CascadeMux I__4464 (
            .O(N__29199),
            .I(N__29196));
    InMux I__4463 (
            .O(N__29196),
            .I(N__29193));
    LocalMux I__4462 (
            .O(N__29193),
            .I(N__29190));
    Span4Mux_h I__4461 (
            .O(N__29190),
            .I(N__29186));
    InMux I__4460 (
            .O(N__29189),
            .I(N__29182));
    Span4Mux_v I__4459 (
            .O(N__29186),
            .I(N__29179));
    InMux I__4458 (
            .O(N__29185),
            .I(N__29176));
    LocalMux I__4457 (
            .O(N__29182),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__4456 (
            .O(N__29179),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__4455 (
            .O(N__29176),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__4454 (
            .O(N__29169),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__4453 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__4452 (
            .O(N__29163),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    CascadeMux I__4451 (
            .O(N__29160),
            .I(N__29156));
    InMux I__4450 (
            .O(N__29159),
            .I(N__29153));
    InMux I__4449 (
            .O(N__29156),
            .I(N__29150));
    LocalMux I__4448 (
            .O(N__29153),
            .I(N__29147));
    LocalMux I__4447 (
            .O(N__29150),
            .I(N__29144));
    Span4Mux_v I__4446 (
            .O(N__29147),
            .I(N__29140));
    Span4Mux_h I__4445 (
            .O(N__29144),
            .I(N__29137));
    InMux I__4444 (
            .O(N__29143),
            .I(N__29134));
    Odrv4 I__4443 (
            .O(N__29140),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv4 I__4442 (
            .O(N__29137),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__4441 (
            .O(N__29134),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__4440 (
            .O(N__29127),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__4439 (
            .O(N__29124),
            .I(N__29121));
    LocalMux I__4438 (
            .O(N__29121),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__4437 (
            .O(N__29118),
            .I(N__29115));
    LocalMux I__4436 (
            .O(N__29115),
            .I(N__29110));
    InMux I__4435 (
            .O(N__29114),
            .I(N__29105));
    InMux I__4434 (
            .O(N__29113),
            .I(N__29105));
    Span4Mux_v I__4433 (
            .O(N__29110),
            .I(N__29100));
    LocalMux I__4432 (
            .O(N__29105),
            .I(N__29100));
    Odrv4 I__4431 (
            .O(N__29100),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__4430 (
            .O(N__29097),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__4429 (
            .O(N__29094),
            .I(N__29091));
    LocalMux I__4428 (
            .O(N__29091),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__4427 (
            .O(N__29088),
            .I(N__29084));
    CascadeMux I__4426 (
            .O(N__29087),
            .I(N__29080));
    LocalMux I__4425 (
            .O(N__29084),
            .I(N__29077));
    InMux I__4424 (
            .O(N__29083),
            .I(N__29074));
    InMux I__4423 (
            .O(N__29080),
            .I(N__29071));
    Span4Mux_v I__4422 (
            .O(N__29077),
            .I(N__29066));
    LocalMux I__4421 (
            .O(N__29074),
            .I(N__29066));
    LocalMux I__4420 (
            .O(N__29071),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__4419 (
            .O(N__29066),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__4418 (
            .O(N__29061),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__4417 (
            .O(N__29058),
            .I(N__29055));
    LocalMux I__4416 (
            .O(N__29055),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__4415 (
            .O(N__29052),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__4414 (
            .O(N__29049),
            .I(N__29046));
    LocalMux I__4413 (
            .O(N__29046),
            .I(\phase_controller_inst1.stoper_hc.un4_start_0 ));
    InMux I__4412 (
            .O(N__29043),
            .I(N__29034));
    InMux I__4411 (
            .O(N__29042),
            .I(N__29034));
    InMux I__4410 (
            .O(N__29041),
            .I(N__29034));
    LocalMux I__4409 (
            .O(N__29034),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__4408 (
            .O(N__29031),
            .I(N__29028));
    LocalMux I__4407 (
            .O(N__29028),
            .I(N__29025));
    Odrv12 I__4406 (
            .O(N__29025),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__4405 (
            .O(N__29022),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__4404 (
            .O(N__29019),
            .I(N__29016));
    LocalMux I__4403 (
            .O(N__29016),
            .I(N__29013));
    Span4Mux_v I__4402 (
            .O(N__29013),
            .I(N__29009));
    InMux I__4401 (
            .O(N__29012),
            .I(N__29006));
    Span4Mux_v I__4400 (
            .O(N__29009),
            .I(N__29001));
    LocalMux I__4399 (
            .O(N__29006),
            .I(N__29001));
    Span4Mux_v I__4398 (
            .O(N__29001),
            .I(N__28998));
    Odrv4 I__4397 (
            .O(N__28998),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__4396 (
            .O(N__28995),
            .I(N__28992));
    LocalMux I__4395 (
            .O(N__28992),
            .I(N__28989));
    Span4Mux_v I__4394 (
            .O(N__28989),
            .I(N__28985));
    InMux I__4393 (
            .O(N__28988),
            .I(N__28982));
    Sp12to4 I__4392 (
            .O(N__28985),
            .I(N__28978));
    LocalMux I__4391 (
            .O(N__28982),
            .I(N__28975));
    InMux I__4390 (
            .O(N__28981),
            .I(N__28972));
    Span12Mux_h I__4389 (
            .O(N__28978),
            .I(N__28967));
    Span12Mux_v I__4388 (
            .O(N__28975),
            .I(N__28967));
    LocalMux I__4387 (
            .O(N__28972),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv12 I__4386 (
            .O(N__28967),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__4385 (
            .O(N__28962),
            .I(N__28959));
    LocalMux I__4384 (
            .O(N__28959),
            .I(N__28940));
    InMux I__4383 (
            .O(N__28958),
            .I(N__28931));
    InMux I__4382 (
            .O(N__28957),
            .I(N__28931));
    InMux I__4381 (
            .O(N__28956),
            .I(N__28931));
    InMux I__4380 (
            .O(N__28955),
            .I(N__28931));
    InMux I__4379 (
            .O(N__28954),
            .I(N__28924));
    InMux I__4378 (
            .O(N__28953),
            .I(N__28924));
    InMux I__4377 (
            .O(N__28952),
            .I(N__28924));
    InMux I__4376 (
            .O(N__28951),
            .I(N__28911));
    InMux I__4375 (
            .O(N__28950),
            .I(N__28911));
    InMux I__4374 (
            .O(N__28949),
            .I(N__28911));
    InMux I__4373 (
            .O(N__28948),
            .I(N__28911));
    InMux I__4372 (
            .O(N__28947),
            .I(N__28911));
    InMux I__4371 (
            .O(N__28946),
            .I(N__28911));
    InMux I__4370 (
            .O(N__28945),
            .I(N__28901));
    InMux I__4369 (
            .O(N__28944),
            .I(N__28901));
    InMux I__4368 (
            .O(N__28943),
            .I(N__28901));
    Span4Mux_h I__4367 (
            .O(N__28940),
            .I(N__28894));
    LocalMux I__4366 (
            .O(N__28931),
            .I(N__28894));
    LocalMux I__4365 (
            .O(N__28924),
            .I(N__28894));
    LocalMux I__4364 (
            .O(N__28911),
            .I(N__28891));
    InMux I__4363 (
            .O(N__28910),
            .I(N__28884));
    InMux I__4362 (
            .O(N__28909),
            .I(N__28884));
    InMux I__4361 (
            .O(N__28908),
            .I(N__28884));
    LocalMux I__4360 (
            .O(N__28901),
            .I(N__28877));
    Span4Mux_v I__4359 (
            .O(N__28894),
            .I(N__28873));
    Span4Mux_h I__4358 (
            .O(N__28891),
            .I(N__28868));
    LocalMux I__4357 (
            .O(N__28884),
            .I(N__28868));
    InMux I__4356 (
            .O(N__28883),
            .I(N__28863));
    InMux I__4355 (
            .O(N__28882),
            .I(N__28863));
    InMux I__4354 (
            .O(N__28881),
            .I(N__28858));
    InMux I__4353 (
            .O(N__28880),
            .I(N__28858));
    Span4Mux_h I__4352 (
            .O(N__28877),
            .I(N__28855));
    InMux I__4351 (
            .O(N__28876),
            .I(N__28852));
    Odrv4 I__4350 (
            .O(N__28873),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__4349 (
            .O(N__28868),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__4348 (
            .O(N__28863),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__4347 (
            .O(N__28858),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__4346 (
            .O(N__28855),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__4345 (
            .O(N__28852),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__4344 (
            .O(N__28839),
            .I(N__28836));
    LocalMux I__4343 (
            .O(N__28836),
            .I(N__28833));
    Span4Mux_v I__4342 (
            .O(N__28833),
            .I(N__28829));
    CascadeMux I__4341 (
            .O(N__28832),
            .I(N__28825));
    Span4Mux_v I__4340 (
            .O(N__28829),
            .I(N__28822));
    InMux I__4339 (
            .O(N__28828),
            .I(N__28819));
    InMux I__4338 (
            .O(N__28825),
            .I(N__28816));
    Odrv4 I__4337 (
            .O(N__28822),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__4336 (
            .O(N__28819),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__4335 (
            .O(N__28816),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__4334 (
            .O(N__28809),
            .I(N__28806));
    LocalMux I__4333 (
            .O(N__28806),
            .I(N__28803));
    Span4Mux_h I__4332 (
            .O(N__28803),
            .I(N__28797));
    InMux I__4331 (
            .O(N__28802),
            .I(N__28794));
    InMux I__4330 (
            .O(N__28801),
            .I(N__28789));
    InMux I__4329 (
            .O(N__28800),
            .I(N__28789));
    Odrv4 I__4328 (
            .O(N__28797),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__4327 (
            .O(N__28794),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__4326 (
            .O(N__28789),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__4325 (
            .O(N__28782),
            .I(N__28779));
    InMux I__4324 (
            .O(N__28779),
            .I(N__28773));
    InMux I__4323 (
            .O(N__28778),
            .I(N__28770));
    InMux I__4322 (
            .O(N__28777),
            .I(N__28767));
    InMux I__4321 (
            .O(N__28776),
            .I(N__28762));
    LocalMux I__4320 (
            .O(N__28773),
            .I(N__28757));
    LocalMux I__4319 (
            .O(N__28770),
            .I(N__28757));
    LocalMux I__4318 (
            .O(N__28767),
            .I(N__28754));
    InMux I__4317 (
            .O(N__28766),
            .I(N__28751));
    InMux I__4316 (
            .O(N__28765),
            .I(N__28748));
    LocalMux I__4315 (
            .O(N__28762),
            .I(N__28745));
    Span4Mux_v I__4314 (
            .O(N__28757),
            .I(N__28740));
    Span4Mux_v I__4313 (
            .O(N__28754),
            .I(N__28740));
    LocalMux I__4312 (
            .O(N__28751),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__4311 (
            .O(N__28748),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv12 I__4310 (
            .O(N__28745),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__4309 (
            .O(N__28740),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__4308 (
            .O(N__28731),
            .I(N__28727));
    InMux I__4307 (
            .O(N__28730),
            .I(N__28724));
    LocalMux I__4306 (
            .O(N__28727),
            .I(N__28721));
    LocalMux I__4305 (
            .O(N__28724),
            .I(N__28717));
    Span4Mux_h I__4304 (
            .O(N__28721),
            .I(N__28714));
    InMux I__4303 (
            .O(N__28720),
            .I(N__28711));
    Odrv12 I__4302 (
            .O(N__28717),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    Odrv4 I__4301 (
            .O(N__28714),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    LocalMux I__4300 (
            .O(N__28711),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    InMux I__4299 (
            .O(N__28704),
            .I(N__28700));
    CascadeMux I__4298 (
            .O(N__28703),
            .I(N__28697));
    LocalMux I__4297 (
            .O(N__28700),
            .I(N__28694));
    InMux I__4296 (
            .O(N__28697),
            .I(N__28691));
    Span4Mux_v I__4295 (
            .O(N__28694),
            .I(N__28688));
    LocalMux I__4294 (
            .O(N__28691),
            .I(N__28685));
    Odrv4 I__4293 (
            .O(N__28688),
            .I(\phase_controller_inst2.stoper_tr.counter ));
    Odrv4 I__4292 (
            .O(N__28685),
            .I(\phase_controller_inst2.stoper_tr.counter ));
    InMux I__4291 (
            .O(N__28680),
            .I(N__28675));
    InMux I__4290 (
            .O(N__28679),
            .I(N__28670));
    InMux I__4289 (
            .O(N__28678),
            .I(N__28670));
    LocalMux I__4288 (
            .O(N__28675),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ));
    LocalMux I__4287 (
            .O(N__28670),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ));
    InMux I__4286 (
            .O(N__28665),
            .I(N__28660));
    InMux I__4285 (
            .O(N__28664),
            .I(N__28655));
    InMux I__4284 (
            .O(N__28663),
            .I(N__28655));
    LocalMux I__4283 (
            .O(N__28660),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ));
    LocalMux I__4282 (
            .O(N__28655),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ));
    InMux I__4281 (
            .O(N__28650),
            .I(N__28647));
    LocalMux I__4280 (
            .O(N__28647),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt24 ));
    CascadeMux I__4279 (
            .O(N__28644),
            .I(N__28641));
    InMux I__4278 (
            .O(N__28641),
            .I(N__28638));
    LocalMux I__4277 (
            .O(N__28638),
            .I(N__28635));
    Odrv4 I__4276 (
            .O(N__28635),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt16 ));
    InMux I__4275 (
            .O(N__28632),
            .I(N__28625));
    InMux I__4274 (
            .O(N__28631),
            .I(N__28625));
    InMux I__4273 (
            .O(N__28630),
            .I(N__28622));
    LocalMux I__4272 (
            .O(N__28625),
            .I(N__28619));
    LocalMux I__4271 (
            .O(N__28622),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ));
    Odrv4 I__4270 (
            .O(N__28619),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ));
    CascadeMux I__4269 (
            .O(N__28614),
            .I(N__28610));
    CascadeMux I__4268 (
            .O(N__28613),
            .I(N__28607));
    InMux I__4267 (
            .O(N__28610),
            .I(N__28601));
    InMux I__4266 (
            .O(N__28607),
            .I(N__28601));
    InMux I__4265 (
            .O(N__28606),
            .I(N__28598));
    LocalMux I__4264 (
            .O(N__28601),
            .I(N__28595));
    LocalMux I__4263 (
            .O(N__28598),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ));
    Odrv4 I__4262 (
            .O(N__28595),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ));
    InMux I__4261 (
            .O(N__28590),
            .I(N__28587));
    LocalMux I__4260 (
            .O(N__28587),
            .I(N__28584));
    Odrv4 I__4259 (
            .O(N__28584),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ));
    InMux I__4258 (
            .O(N__28581),
            .I(N__28578));
    LocalMux I__4257 (
            .O(N__28578),
            .I(N__28575));
    Span4Mux_h I__4256 (
            .O(N__28575),
            .I(N__28572));
    Odrv4 I__4255 (
            .O(N__28572),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ));
    InMux I__4254 (
            .O(N__28569),
            .I(N__28566));
    LocalMux I__4253 (
            .O(N__28566),
            .I(N__28563));
    Odrv12 I__4252 (
            .O(N__28563),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__4251 (
            .O(N__28560),
            .I(N__28553));
    InMux I__4250 (
            .O(N__28559),
            .I(N__28553));
    InMux I__4249 (
            .O(N__28558),
            .I(N__28550));
    LocalMux I__4248 (
            .O(N__28553),
            .I(N__28547));
    LocalMux I__4247 (
            .O(N__28550),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ));
    Odrv4 I__4246 (
            .O(N__28547),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ));
    InMux I__4245 (
            .O(N__28542),
            .I(N__28535));
    InMux I__4244 (
            .O(N__28541),
            .I(N__28535));
    InMux I__4243 (
            .O(N__28540),
            .I(N__28532));
    LocalMux I__4242 (
            .O(N__28535),
            .I(N__28529));
    LocalMux I__4241 (
            .O(N__28532),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ));
    Odrv4 I__4240 (
            .O(N__28529),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ));
    CascadeMux I__4239 (
            .O(N__28524),
            .I(N__28521));
    InMux I__4238 (
            .O(N__28521),
            .I(N__28518));
    LocalMux I__4237 (
            .O(N__28518),
            .I(N__28515));
    Span4Mux_h I__4236 (
            .O(N__28515),
            .I(N__28512));
    Odrv4 I__4235 (
            .O(N__28512),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt18 ));
    InMux I__4234 (
            .O(N__28509),
            .I(N__28506));
    LocalMux I__4233 (
            .O(N__28506),
            .I(N__28503));
    Odrv4 I__4232 (
            .O(N__28503),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ));
    CascadeMux I__4231 (
            .O(N__28500),
            .I(N__28497));
    InMux I__4230 (
            .O(N__28497),
            .I(N__28494));
    LocalMux I__4229 (
            .O(N__28494),
            .I(N__28491));
    Span4Mux_h I__4228 (
            .O(N__28491),
            .I(N__28488));
    Odrv4 I__4227 (
            .O(N__28488),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ));
    CascadeMux I__4226 (
            .O(N__28485),
            .I(N__28482));
    InMux I__4225 (
            .O(N__28482),
            .I(N__28479));
    LocalMux I__4224 (
            .O(N__28479),
            .I(N__28476));
    Odrv4 I__4223 (
            .O(N__28476),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ));
    InMux I__4222 (
            .O(N__28473),
            .I(bfn_11_10_0_));
    InMux I__4221 (
            .O(N__28470),
            .I(N__28465));
    InMux I__4220 (
            .O(N__28469),
            .I(N__28462));
    InMux I__4219 (
            .O(N__28468),
            .I(N__28459));
    LocalMux I__4218 (
            .O(N__28465),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    LocalMux I__4217 (
            .O(N__28462),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    LocalMux I__4216 (
            .O(N__28459),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    InMux I__4215 (
            .O(N__28452),
            .I(N__28447));
    InMux I__4214 (
            .O(N__28451),
            .I(N__28444));
    InMux I__4213 (
            .O(N__28450),
            .I(N__28441));
    LocalMux I__4212 (
            .O(N__28447),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    LocalMux I__4211 (
            .O(N__28444),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    LocalMux I__4210 (
            .O(N__28441),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    InMux I__4209 (
            .O(N__28434),
            .I(N__28431));
    LocalMux I__4208 (
            .O(N__28431),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt30 ));
    CascadeMux I__4207 (
            .O(N__28428),
            .I(N__28425));
    InMux I__4206 (
            .O(N__28425),
            .I(N__28422));
    LocalMux I__4205 (
            .O(N__28422),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ));
    InMux I__4204 (
            .O(N__28419),
            .I(N__28413));
    InMux I__4203 (
            .O(N__28418),
            .I(N__28408));
    InMux I__4202 (
            .O(N__28417),
            .I(N__28408));
    InMux I__4201 (
            .O(N__28416),
            .I(N__28405));
    LocalMux I__4200 (
            .O(N__28413),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ));
    LocalMux I__4199 (
            .O(N__28408),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ));
    LocalMux I__4198 (
            .O(N__28405),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ));
    InMux I__4197 (
            .O(N__28398),
            .I(N__28393));
    InMux I__4196 (
            .O(N__28397),
            .I(N__28390));
    InMux I__4195 (
            .O(N__28396),
            .I(N__28387));
    LocalMux I__4194 (
            .O(N__28393),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    LocalMux I__4193 (
            .O(N__28390),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    LocalMux I__4192 (
            .O(N__28387),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    InMux I__4191 (
            .O(N__28380),
            .I(N__28375));
    InMux I__4190 (
            .O(N__28379),
            .I(N__28372));
    InMux I__4189 (
            .O(N__28378),
            .I(N__28369));
    LocalMux I__4188 (
            .O(N__28375),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    LocalMux I__4187 (
            .O(N__28372),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    LocalMux I__4186 (
            .O(N__28369),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    InMux I__4185 (
            .O(N__28362),
            .I(N__28359));
    LocalMux I__4184 (
            .O(N__28359),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt28 ));
    InMux I__4183 (
            .O(N__28356),
            .I(N__28352));
    InMux I__4182 (
            .O(N__28355),
            .I(N__28349));
    LocalMux I__4181 (
            .O(N__28352),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ));
    LocalMux I__4180 (
            .O(N__28349),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ));
    CascadeMux I__4179 (
            .O(N__28344),
            .I(N__28341));
    InMux I__4178 (
            .O(N__28341),
            .I(N__28338));
    LocalMux I__4177 (
            .O(N__28338),
            .I(\phase_controller_inst2.stoper_tr.counter_i_11 ));
    InMux I__4176 (
            .O(N__28335),
            .I(N__28331));
    InMux I__4175 (
            .O(N__28334),
            .I(N__28328));
    LocalMux I__4174 (
            .O(N__28331),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ));
    LocalMux I__4173 (
            .O(N__28328),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ));
    CascadeMux I__4172 (
            .O(N__28323),
            .I(N__28320));
    InMux I__4171 (
            .O(N__28320),
            .I(N__28317));
    LocalMux I__4170 (
            .O(N__28317),
            .I(\phase_controller_inst2.stoper_tr.counter_i_12 ));
    InMux I__4169 (
            .O(N__28314),
            .I(N__28310));
    InMux I__4168 (
            .O(N__28313),
            .I(N__28307));
    LocalMux I__4167 (
            .O(N__28310),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ));
    LocalMux I__4166 (
            .O(N__28307),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ));
    CascadeMux I__4165 (
            .O(N__28302),
            .I(N__28299));
    InMux I__4164 (
            .O(N__28299),
            .I(N__28296));
    LocalMux I__4163 (
            .O(N__28296),
            .I(\phase_controller_inst2.stoper_tr.counter_i_13 ));
    InMux I__4162 (
            .O(N__28293),
            .I(N__28289));
    InMux I__4161 (
            .O(N__28292),
            .I(N__28286));
    LocalMux I__4160 (
            .O(N__28289),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ));
    LocalMux I__4159 (
            .O(N__28286),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ));
    CascadeMux I__4158 (
            .O(N__28281),
            .I(N__28278));
    InMux I__4157 (
            .O(N__28278),
            .I(N__28275));
    LocalMux I__4156 (
            .O(N__28275),
            .I(\phase_controller_inst2.stoper_tr.counter_i_14 ));
    InMux I__4155 (
            .O(N__28272),
            .I(N__28268));
    InMux I__4154 (
            .O(N__28271),
            .I(N__28265));
    LocalMux I__4153 (
            .O(N__28268),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ));
    LocalMux I__4152 (
            .O(N__28265),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ));
    CascadeMux I__4151 (
            .O(N__28260),
            .I(N__28257));
    InMux I__4150 (
            .O(N__28257),
            .I(N__28254));
    LocalMux I__4149 (
            .O(N__28254),
            .I(\phase_controller_inst2.stoper_tr.counter_i_15 ));
    InMux I__4148 (
            .O(N__28251),
            .I(N__28247));
    InMux I__4147 (
            .O(N__28250),
            .I(N__28244));
    LocalMux I__4146 (
            .O(N__28247),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ));
    LocalMux I__4145 (
            .O(N__28244),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ));
    CascadeMux I__4144 (
            .O(N__28239),
            .I(N__28236));
    InMux I__4143 (
            .O(N__28236),
            .I(N__28233));
    LocalMux I__4142 (
            .O(N__28233),
            .I(\phase_controller_inst2.stoper_tr.counter_i_3 ));
    InMux I__4141 (
            .O(N__28230),
            .I(N__28226));
    InMux I__4140 (
            .O(N__28229),
            .I(N__28223));
    LocalMux I__4139 (
            .O(N__28226),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ));
    LocalMux I__4138 (
            .O(N__28223),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ));
    CascadeMux I__4137 (
            .O(N__28218),
            .I(N__28215));
    InMux I__4136 (
            .O(N__28215),
            .I(N__28212));
    LocalMux I__4135 (
            .O(N__28212),
            .I(\phase_controller_inst2.stoper_tr.counter_i_4 ));
    InMux I__4134 (
            .O(N__28209),
            .I(N__28205));
    InMux I__4133 (
            .O(N__28208),
            .I(N__28202));
    LocalMux I__4132 (
            .O(N__28205),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ));
    LocalMux I__4131 (
            .O(N__28202),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ));
    CascadeMux I__4130 (
            .O(N__28197),
            .I(N__28194));
    InMux I__4129 (
            .O(N__28194),
            .I(N__28191));
    LocalMux I__4128 (
            .O(N__28191),
            .I(\phase_controller_inst2.stoper_tr.counter_i_5 ));
    InMux I__4127 (
            .O(N__28188),
            .I(N__28184));
    InMux I__4126 (
            .O(N__28187),
            .I(N__28181));
    LocalMux I__4125 (
            .O(N__28184),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ));
    LocalMux I__4124 (
            .O(N__28181),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ));
    CascadeMux I__4123 (
            .O(N__28176),
            .I(N__28173));
    InMux I__4122 (
            .O(N__28173),
            .I(N__28170));
    LocalMux I__4121 (
            .O(N__28170),
            .I(\phase_controller_inst2.stoper_tr.counter_i_6 ));
    InMux I__4120 (
            .O(N__28167),
            .I(N__28163));
    InMux I__4119 (
            .O(N__28166),
            .I(N__28160));
    LocalMux I__4118 (
            .O(N__28163),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ));
    LocalMux I__4117 (
            .O(N__28160),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ));
    CascadeMux I__4116 (
            .O(N__28155),
            .I(N__28152));
    InMux I__4115 (
            .O(N__28152),
            .I(N__28149));
    LocalMux I__4114 (
            .O(N__28149),
            .I(\phase_controller_inst2.stoper_tr.counter_i_7 ));
    InMux I__4113 (
            .O(N__28146),
            .I(N__28142));
    InMux I__4112 (
            .O(N__28145),
            .I(N__28139));
    LocalMux I__4111 (
            .O(N__28142),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ));
    LocalMux I__4110 (
            .O(N__28139),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ));
    CascadeMux I__4109 (
            .O(N__28134),
            .I(N__28131));
    InMux I__4108 (
            .O(N__28131),
            .I(N__28128));
    LocalMux I__4107 (
            .O(N__28128),
            .I(\phase_controller_inst2.stoper_tr.counter_i_8 ));
    InMux I__4106 (
            .O(N__28125),
            .I(N__28121));
    InMux I__4105 (
            .O(N__28124),
            .I(N__28118));
    LocalMux I__4104 (
            .O(N__28121),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ));
    LocalMux I__4103 (
            .O(N__28118),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ));
    CascadeMux I__4102 (
            .O(N__28113),
            .I(N__28110));
    InMux I__4101 (
            .O(N__28110),
            .I(N__28107));
    LocalMux I__4100 (
            .O(N__28107),
            .I(\phase_controller_inst2.stoper_tr.counter_i_9 ));
    InMux I__4099 (
            .O(N__28104),
            .I(N__28100));
    InMux I__4098 (
            .O(N__28103),
            .I(N__28097));
    LocalMux I__4097 (
            .O(N__28100),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ));
    LocalMux I__4096 (
            .O(N__28097),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ));
    CascadeMux I__4095 (
            .O(N__28092),
            .I(N__28089));
    InMux I__4094 (
            .O(N__28089),
            .I(N__28086));
    LocalMux I__4093 (
            .O(N__28086),
            .I(\phase_controller_inst2.stoper_tr.counter_i_10 ));
    IoInMux I__4092 (
            .O(N__28083),
            .I(N__28080));
    LocalMux I__4091 (
            .O(N__28080),
            .I(N__28077));
    Span4Mux_s1_v I__4090 (
            .O(N__28077),
            .I(N__28074));
    Odrv4 I__4089 (
            .O(N__28074),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    CascadeMux I__4088 (
            .O(N__28071),
            .I(N__28068));
    InMux I__4087 (
            .O(N__28068),
            .I(N__28065));
    LocalMux I__4086 (
            .O(N__28065),
            .I(\phase_controller_inst2.stoper_hc.un4_start_0 ));
    InMux I__4085 (
            .O(N__28062),
            .I(N__28056));
    InMux I__4084 (
            .O(N__28061),
            .I(N__28056));
    LocalMux I__4083 (
            .O(N__28056),
            .I(N__28052));
    InMux I__4082 (
            .O(N__28055),
            .I(N__28048));
    Span4Mux_v I__4081 (
            .O(N__28052),
            .I(N__28045));
    InMux I__4080 (
            .O(N__28051),
            .I(N__28042));
    LocalMux I__4079 (
            .O(N__28048),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__4078 (
            .O(N__28045),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__4077 (
            .O(N__28042),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__4076 (
            .O(N__28035),
            .I(N__28030));
    InMux I__4075 (
            .O(N__28034),
            .I(N__28024));
    InMux I__4074 (
            .O(N__28033),
            .I(N__28021));
    LocalMux I__4073 (
            .O(N__28030),
            .I(N__28018));
    InMux I__4072 (
            .O(N__28029),
            .I(N__28015));
    InMux I__4071 (
            .O(N__28028),
            .I(N__28012));
    InMux I__4070 (
            .O(N__28027),
            .I(N__28009));
    LocalMux I__4069 (
            .O(N__28024),
            .I(N__28006));
    LocalMux I__4068 (
            .O(N__28021),
            .I(N__27999));
    Span4Mux_v I__4067 (
            .O(N__28018),
            .I(N__27999));
    LocalMux I__4066 (
            .O(N__28015),
            .I(N__27999));
    LocalMux I__4065 (
            .O(N__28012),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__4064 (
            .O(N__28009),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__4063 (
            .O(N__28006),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__4062 (
            .O(N__27999),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__4061 (
            .O(N__27990),
            .I(N__27986));
    InMux I__4060 (
            .O(N__27989),
            .I(N__27982));
    LocalMux I__4059 (
            .O(N__27986),
            .I(N__27979));
    InMux I__4058 (
            .O(N__27985),
            .I(N__27976));
    LocalMux I__4057 (
            .O(N__27982),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    Odrv4 I__4056 (
            .O(N__27979),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__4055 (
            .O(N__27976),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__4054 (
            .O(N__27969),
            .I(N__27965));
    InMux I__4053 (
            .O(N__27968),
            .I(N__27962));
    LocalMux I__4052 (
            .O(N__27965),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ));
    LocalMux I__4051 (
            .O(N__27962),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ));
    CascadeMux I__4050 (
            .O(N__27957),
            .I(N__27954));
    InMux I__4049 (
            .O(N__27954),
            .I(N__27951));
    LocalMux I__4048 (
            .O(N__27951),
            .I(\phase_controller_inst2.stoper_tr.counter_i_0 ));
    InMux I__4047 (
            .O(N__27948),
            .I(N__27944));
    InMux I__4046 (
            .O(N__27947),
            .I(N__27941));
    LocalMux I__4045 (
            .O(N__27944),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ));
    LocalMux I__4044 (
            .O(N__27941),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ));
    CascadeMux I__4043 (
            .O(N__27936),
            .I(N__27933));
    InMux I__4042 (
            .O(N__27933),
            .I(N__27930));
    LocalMux I__4041 (
            .O(N__27930),
            .I(\phase_controller_inst2.stoper_tr.counter_i_1 ));
    InMux I__4040 (
            .O(N__27927),
            .I(N__27923));
    InMux I__4039 (
            .O(N__27926),
            .I(N__27920));
    LocalMux I__4038 (
            .O(N__27923),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ));
    LocalMux I__4037 (
            .O(N__27920),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ));
    CascadeMux I__4036 (
            .O(N__27915),
            .I(N__27912));
    InMux I__4035 (
            .O(N__27912),
            .I(N__27909));
    LocalMux I__4034 (
            .O(N__27909),
            .I(\phase_controller_inst2.stoper_tr.counter_i_2 ));
    CascadeMux I__4033 (
            .O(N__27906),
            .I(N__27902));
    InMux I__4032 (
            .O(N__27905),
            .I(N__27898));
    InMux I__4031 (
            .O(N__27902),
            .I(N__27895));
    InMux I__4030 (
            .O(N__27901),
            .I(N__27892));
    LocalMux I__4029 (
            .O(N__27898),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    LocalMux I__4028 (
            .O(N__27895),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    LocalMux I__4027 (
            .O(N__27892),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__4026 (
            .O(N__27885),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__4025 (
            .O(N__27882),
            .I(N__27878));
    InMux I__4024 (
            .O(N__27881),
            .I(N__27874));
    InMux I__4023 (
            .O(N__27878),
            .I(N__27871));
    InMux I__4022 (
            .O(N__27877),
            .I(N__27868));
    LocalMux I__4021 (
            .O(N__27874),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__4020 (
            .O(N__27871),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__4019 (
            .O(N__27868),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__4018 (
            .O(N__27861),
            .I(bfn_10_23_0_));
    CascadeMux I__4017 (
            .O(N__27858),
            .I(N__27854));
    InMux I__4016 (
            .O(N__27857),
            .I(N__27850));
    InMux I__4015 (
            .O(N__27854),
            .I(N__27847));
    InMux I__4014 (
            .O(N__27853),
            .I(N__27844));
    LocalMux I__4013 (
            .O(N__27850),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__4012 (
            .O(N__27847),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__4011 (
            .O(N__27844),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__4010 (
            .O(N__27837),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__4009 (
            .O(N__27834),
            .I(N__27830));
    InMux I__4008 (
            .O(N__27833),
            .I(N__27827));
    LocalMux I__4007 (
            .O(N__27830),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    LocalMux I__4006 (
            .O(N__27827),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    CascadeMux I__4005 (
            .O(N__27822),
            .I(N__27818));
    InMux I__4004 (
            .O(N__27821),
            .I(N__27814));
    InMux I__4003 (
            .O(N__27818),
            .I(N__27811));
    InMux I__4002 (
            .O(N__27817),
            .I(N__27808));
    LocalMux I__4001 (
            .O(N__27814),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    LocalMux I__4000 (
            .O(N__27811),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    LocalMux I__3999 (
            .O(N__27808),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__3998 (
            .O(N__27801),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__3997 (
            .O(N__27798),
            .I(N__27794));
    InMux I__3996 (
            .O(N__27797),
            .I(N__27791));
    LocalMux I__3995 (
            .O(N__27794),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    LocalMux I__3994 (
            .O(N__27791),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CascadeMux I__3993 (
            .O(N__27786),
            .I(N__27782));
    InMux I__3992 (
            .O(N__27785),
            .I(N__27778));
    InMux I__3991 (
            .O(N__27782),
            .I(N__27775));
    InMux I__3990 (
            .O(N__27781),
            .I(N__27772));
    LocalMux I__3989 (
            .O(N__27778),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    LocalMux I__3988 (
            .O(N__27775),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    LocalMux I__3987 (
            .O(N__27772),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__3986 (
            .O(N__27765),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__3985 (
            .O(N__27762),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__3984 (
            .O(N__27759),
            .I(N__27755));
    InMux I__3983 (
            .O(N__27758),
            .I(N__27751));
    InMux I__3982 (
            .O(N__27755),
            .I(N__27748));
    InMux I__3981 (
            .O(N__27754),
            .I(N__27745));
    LocalMux I__3980 (
            .O(N__27751),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    LocalMux I__3979 (
            .O(N__27748),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    LocalMux I__3978 (
            .O(N__27745),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__3977 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__3976 (
            .O(N__27735),
            .I(N__27730));
    InMux I__3975 (
            .O(N__27734),
            .I(N__27727));
    CascadeMux I__3974 (
            .O(N__27733),
            .I(N__27724));
    Span4Mux_v I__3973 (
            .O(N__27730),
            .I(N__27718));
    LocalMux I__3972 (
            .O(N__27727),
            .I(N__27718));
    InMux I__3971 (
            .O(N__27724),
            .I(N__27713));
    InMux I__3970 (
            .O(N__27723),
            .I(N__27713));
    Span4Mux_v I__3969 (
            .O(N__27718),
            .I(N__27710));
    LocalMux I__3968 (
            .O(N__27713),
            .I(N__27707));
    Odrv4 I__3967 (
            .O(N__27710),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv12 I__3966 (
            .O(N__27707),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__3965 (
            .O(N__27702),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__3964 (
            .O(N__27699),
            .I(N__27695));
    InMux I__3963 (
            .O(N__27698),
            .I(N__27691));
    InMux I__3962 (
            .O(N__27695),
            .I(N__27688));
    InMux I__3961 (
            .O(N__27694),
            .I(N__27685));
    LocalMux I__3960 (
            .O(N__27691),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__3959 (
            .O(N__27688),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__3958 (
            .O(N__27685),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__3957 (
            .O(N__27678),
            .I(N__27674));
    InMux I__3956 (
            .O(N__27677),
            .I(N__27669));
    LocalMux I__3955 (
            .O(N__27674),
            .I(N__27666));
    InMux I__3954 (
            .O(N__27673),
            .I(N__27663));
    InMux I__3953 (
            .O(N__27672),
            .I(N__27660));
    LocalMux I__3952 (
            .O(N__27669),
            .I(N__27657));
    Span4Mux_v I__3951 (
            .O(N__27666),
            .I(N__27652));
    LocalMux I__3950 (
            .O(N__27663),
            .I(N__27652));
    LocalMux I__3949 (
            .O(N__27660),
            .I(N__27649));
    Span4Mux_h I__3948 (
            .O(N__27657),
            .I(N__27646));
    Span4Mux_v I__3947 (
            .O(N__27652),
            .I(N__27641));
    Span4Mux_h I__3946 (
            .O(N__27649),
            .I(N__27641));
    Odrv4 I__3945 (
            .O(N__27646),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__3944 (
            .O(N__27641),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__3943 (
            .O(N__27636),
            .I(bfn_10_22_0_));
    CascadeMux I__3942 (
            .O(N__27633),
            .I(N__27629));
    InMux I__3941 (
            .O(N__27632),
            .I(N__27625));
    InMux I__3940 (
            .O(N__27629),
            .I(N__27622));
    InMux I__3939 (
            .O(N__27628),
            .I(N__27619));
    LocalMux I__3938 (
            .O(N__27625),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    LocalMux I__3937 (
            .O(N__27622),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    LocalMux I__3936 (
            .O(N__27619),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    CascadeMux I__3935 (
            .O(N__27612),
            .I(N__27609));
    InMux I__3934 (
            .O(N__27609),
            .I(N__27605));
    InMux I__3933 (
            .O(N__27608),
            .I(N__27600));
    LocalMux I__3932 (
            .O(N__27605),
            .I(N__27597));
    InMux I__3931 (
            .O(N__27604),
            .I(N__27594));
    InMux I__3930 (
            .O(N__27603),
            .I(N__27591));
    LocalMux I__3929 (
            .O(N__27600),
            .I(N__27588));
    Span4Mux_v I__3928 (
            .O(N__27597),
            .I(N__27581));
    LocalMux I__3927 (
            .O(N__27594),
            .I(N__27581));
    LocalMux I__3926 (
            .O(N__27591),
            .I(N__27581));
    Span4Mux_v I__3925 (
            .O(N__27588),
            .I(N__27578));
    Span4Mux_v I__3924 (
            .O(N__27581),
            .I(N__27575));
    Odrv4 I__3923 (
            .O(N__27578),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__3922 (
            .O(N__27575),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__3921 (
            .O(N__27570),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__3920 (
            .O(N__27567),
            .I(N__27563));
    InMux I__3919 (
            .O(N__27566),
            .I(N__27559));
    InMux I__3918 (
            .O(N__27563),
            .I(N__27556));
    InMux I__3917 (
            .O(N__27562),
            .I(N__27553));
    LocalMux I__3916 (
            .O(N__27559),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    LocalMux I__3915 (
            .O(N__27556),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    LocalMux I__3914 (
            .O(N__27553),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__3913 (
            .O(N__27546),
            .I(N__27542));
    InMux I__3912 (
            .O(N__27545),
            .I(N__27537));
    LocalMux I__3911 (
            .O(N__27542),
            .I(N__27534));
    InMux I__3910 (
            .O(N__27541),
            .I(N__27531));
    InMux I__3909 (
            .O(N__27540),
            .I(N__27528));
    LocalMux I__3908 (
            .O(N__27537),
            .I(N__27523));
    Span4Mux_v I__3907 (
            .O(N__27534),
            .I(N__27523));
    LocalMux I__3906 (
            .O(N__27531),
            .I(N__27518));
    LocalMux I__3905 (
            .O(N__27528),
            .I(N__27518));
    Odrv4 I__3904 (
            .O(N__27523),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv12 I__3903 (
            .O(N__27518),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__3902 (
            .O(N__27513),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__3901 (
            .O(N__27510),
            .I(N__27506));
    InMux I__3900 (
            .O(N__27509),
            .I(N__27502));
    InMux I__3899 (
            .O(N__27506),
            .I(N__27499));
    InMux I__3898 (
            .O(N__27505),
            .I(N__27496));
    LocalMux I__3897 (
            .O(N__27502),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    LocalMux I__3896 (
            .O(N__27499),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    LocalMux I__3895 (
            .O(N__27496),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    CascadeMux I__3894 (
            .O(N__27489),
            .I(N__27486));
    InMux I__3893 (
            .O(N__27486),
            .I(N__27483));
    LocalMux I__3892 (
            .O(N__27483),
            .I(N__27478));
    InMux I__3891 (
            .O(N__27482),
            .I(N__27475));
    InMux I__3890 (
            .O(N__27481),
            .I(N__27471));
    Span4Mux_v I__3889 (
            .O(N__27478),
            .I(N__27466));
    LocalMux I__3888 (
            .O(N__27475),
            .I(N__27466));
    InMux I__3887 (
            .O(N__27474),
            .I(N__27463));
    LocalMux I__3886 (
            .O(N__27471),
            .I(N__27460));
    Sp12to4 I__3885 (
            .O(N__27466),
            .I(N__27455));
    LocalMux I__3884 (
            .O(N__27463),
            .I(N__27455));
    Odrv4 I__3883 (
            .O(N__27460),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv12 I__3882 (
            .O(N__27455),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__3881 (
            .O(N__27450),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__3880 (
            .O(N__27447),
            .I(N__27443));
    InMux I__3879 (
            .O(N__27446),
            .I(N__27439));
    InMux I__3878 (
            .O(N__27443),
            .I(N__27436));
    InMux I__3877 (
            .O(N__27442),
            .I(N__27433));
    LocalMux I__3876 (
            .O(N__27439),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    LocalMux I__3875 (
            .O(N__27436),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    LocalMux I__3874 (
            .O(N__27433),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__3873 (
            .O(N__27426),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__3872 (
            .O(N__27423),
            .I(N__27419));
    InMux I__3871 (
            .O(N__27422),
            .I(N__27415));
    InMux I__3870 (
            .O(N__27419),
            .I(N__27412));
    InMux I__3869 (
            .O(N__27418),
            .I(N__27409));
    LocalMux I__3868 (
            .O(N__27415),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    LocalMux I__3867 (
            .O(N__27412),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    LocalMux I__3866 (
            .O(N__27409),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__3865 (
            .O(N__27402),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__3864 (
            .O(N__27399),
            .I(N__27395));
    InMux I__3863 (
            .O(N__27398),
            .I(N__27391));
    InMux I__3862 (
            .O(N__27395),
            .I(N__27388));
    InMux I__3861 (
            .O(N__27394),
            .I(N__27385));
    LocalMux I__3860 (
            .O(N__27391),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    LocalMux I__3859 (
            .O(N__27388),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    LocalMux I__3858 (
            .O(N__27385),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__3857 (
            .O(N__27378),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__3856 (
            .O(N__27375),
            .I(N__27371));
    InMux I__3855 (
            .O(N__27374),
            .I(N__27367));
    InMux I__3854 (
            .O(N__27371),
            .I(N__27364));
    InMux I__3853 (
            .O(N__27370),
            .I(N__27361));
    LocalMux I__3852 (
            .O(N__27367),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    LocalMux I__3851 (
            .O(N__27364),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    LocalMux I__3850 (
            .O(N__27361),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__3849 (
            .O(N__27354),
            .I(N__27350));
    CascadeMux I__3848 (
            .O(N__27353),
            .I(N__27347));
    LocalMux I__3847 (
            .O(N__27350),
            .I(N__27343));
    InMux I__3846 (
            .O(N__27347),
            .I(N__27340));
    InMux I__3845 (
            .O(N__27346),
            .I(N__27337));
    Span4Mux_v I__3844 (
            .O(N__27343),
            .I(N__27330));
    LocalMux I__3843 (
            .O(N__27340),
            .I(N__27330));
    LocalMux I__3842 (
            .O(N__27337),
            .I(N__27330));
    Span4Mux_v I__3841 (
            .O(N__27330),
            .I(N__27326));
    InMux I__3840 (
            .O(N__27329),
            .I(N__27323));
    Odrv4 I__3839 (
            .O(N__27326),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__3838 (
            .O(N__27323),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__3837 (
            .O(N__27318),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__3836 (
            .O(N__27315),
            .I(N__27311));
    InMux I__3835 (
            .O(N__27314),
            .I(N__27307));
    InMux I__3834 (
            .O(N__27311),
            .I(N__27304));
    InMux I__3833 (
            .O(N__27310),
            .I(N__27301));
    LocalMux I__3832 (
            .O(N__27307),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__3831 (
            .O(N__27304),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__3830 (
            .O(N__27301),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    CascadeMux I__3829 (
            .O(N__27294),
            .I(N__27290));
    InMux I__3828 (
            .O(N__27293),
            .I(N__27286));
    InMux I__3827 (
            .O(N__27290),
            .I(N__27283));
    CascadeMux I__3826 (
            .O(N__27289),
            .I(N__27280));
    LocalMux I__3825 (
            .O(N__27286),
            .I(N__27276));
    LocalMux I__3824 (
            .O(N__27283),
            .I(N__27273));
    InMux I__3823 (
            .O(N__27280),
            .I(N__27270));
    InMux I__3822 (
            .O(N__27279),
            .I(N__27267));
    Span4Mux_v I__3821 (
            .O(N__27276),
            .I(N__27264));
    Sp12to4 I__3820 (
            .O(N__27273),
            .I(N__27257));
    LocalMux I__3819 (
            .O(N__27270),
            .I(N__27257));
    LocalMux I__3818 (
            .O(N__27267),
            .I(N__27257));
    Odrv4 I__3817 (
            .O(N__27264),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv12 I__3816 (
            .O(N__27257),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__3815 (
            .O(N__27252),
            .I(bfn_10_21_0_));
    CascadeMux I__3814 (
            .O(N__27249),
            .I(N__27245));
    InMux I__3813 (
            .O(N__27248),
            .I(N__27241));
    InMux I__3812 (
            .O(N__27245),
            .I(N__27238));
    InMux I__3811 (
            .O(N__27244),
            .I(N__27235));
    LocalMux I__3810 (
            .O(N__27241),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__3809 (
            .O(N__27238),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__3808 (
            .O(N__27235),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    CascadeMux I__3807 (
            .O(N__27228),
            .I(N__27223));
    CascadeMux I__3806 (
            .O(N__27227),
            .I(N__27220));
    InMux I__3805 (
            .O(N__27226),
            .I(N__27217));
    InMux I__3804 (
            .O(N__27223),
            .I(N__27214));
    InMux I__3803 (
            .O(N__27220),
            .I(N__27210));
    LocalMux I__3802 (
            .O(N__27217),
            .I(N__27207));
    LocalMux I__3801 (
            .O(N__27214),
            .I(N__27204));
    InMux I__3800 (
            .O(N__27213),
            .I(N__27201));
    LocalMux I__3799 (
            .O(N__27210),
            .I(N__27198));
    Span4Mux_v I__3798 (
            .O(N__27207),
            .I(N__27195));
    Sp12to4 I__3797 (
            .O(N__27204),
            .I(N__27190));
    LocalMux I__3796 (
            .O(N__27201),
            .I(N__27190));
    Odrv12 I__3795 (
            .O(N__27198),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__3794 (
            .O(N__27195),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv12 I__3793 (
            .O(N__27190),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__3792 (
            .O(N__27183),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__3791 (
            .O(N__27180),
            .I(N__27176));
    InMux I__3790 (
            .O(N__27179),
            .I(N__27172));
    InMux I__3789 (
            .O(N__27176),
            .I(N__27169));
    InMux I__3788 (
            .O(N__27175),
            .I(N__27166));
    LocalMux I__3787 (
            .O(N__27172),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    LocalMux I__3786 (
            .O(N__27169),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    LocalMux I__3785 (
            .O(N__27166),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__3784 (
            .O(N__27159),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__3783 (
            .O(N__27156),
            .I(N__27152));
    InMux I__3782 (
            .O(N__27155),
            .I(N__27148));
    InMux I__3781 (
            .O(N__27152),
            .I(N__27145));
    InMux I__3780 (
            .O(N__27151),
            .I(N__27142));
    LocalMux I__3779 (
            .O(N__27148),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    LocalMux I__3778 (
            .O(N__27145),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    LocalMux I__3777 (
            .O(N__27142),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__3776 (
            .O(N__27135),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__3775 (
            .O(N__27132),
            .I(N__27128));
    InMux I__3774 (
            .O(N__27131),
            .I(N__27124));
    InMux I__3773 (
            .O(N__27128),
            .I(N__27121));
    InMux I__3772 (
            .O(N__27127),
            .I(N__27118));
    LocalMux I__3771 (
            .O(N__27124),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    LocalMux I__3770 (
            .O(N__27121),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    LocalMux I__3769 (
            .O(N__27118),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    CascadeMux I__3768 (
            .O(N__27111),
            .I(N__27107));
    CascadeMux I__3767 (
            .O(N__27110),
            .I(N__27104));
    InMux I__3766 (
            .O(N__27107),
            .I(N__27100));
    InMux I__3765 (
            .O(N__27104),
            .I(N__27095));
    InMux I__3764 (
            .O(N__27103),
            .I(N__27095));
    LocalMux I__3763 (
            .O(N__27100),
            .I(N__27089));
    LocalMux I__3762 (
            .O(N__27095),
            .I(N__27089));
    InMux I__3761 (
            .O(N__27094),
            .I(N__27086));
    Span4Mux_v I__3760 (
            .O(N__27089),
            .I(N__27081));
    LocalMux I__3759 (
            .O(N__27086),
            .I(N__27081));
    Odrv4 I__3758 (
            .O(N__27081),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__3757 (
            .O(N__27078),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__3756 (
            .O(N__27075),
            .I(N__27071));
    InMux I__3755 (
            .O(N__27074),
            .I(N__27067));
    InMux I__3754 (
            .O(N__27071),
            .I(N__27064));
    InMux I__3753 (
            .O(N__27070),
            .I(N__27061));
    LocalMux I__3752 (
            .O(N__27067),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    LocalMux I__3751 (
            .O(N__27064),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    LocalMux I__3750 (
            .O(N__27061),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__3749 (
            .O(N__27054),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__3748 (
            .O(N__27051),
            .I(N__27047));
    InMux I__3747 (
            .O(N__27050),
            .I(N__27043));
    InMux I__3746 (
            .O(N__27047),
            .I(N__27040));
    InMux I__3745 (
            .O(N__27046),
            .I(N__27037));
    LocalMux I__3744 (
            .O(N__27043),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    LocalMux I__3743 (
            .O(N__27040),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    LocalMux I__3742 (
            .O(N__27037),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__3741 (
            .O(N__27030),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__3740 (
            .O(N__27027),
            .I(N__27024));
    LocalMux I__3739 (
            .O(N__27024),
            .I(N__27021));
    Span4Mux_h I__3738 (
            .O(N__27021),
            .I(N__27018));
    Odrv4 I__3737 (
            .O(N__27018),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    CascadeMux I__3736 (
            .O(N__27015),
            .I(N__27011));
    InMux I__3735 (
            .O(N__27014),
            .I(N__27008));
    InMux I__3734 (
            .O(N__27011),
            .I(N__27003));
    LocalMux I__3733 (
            .O(N__27008),
            .I(N__27000));
    InMux I__3732 (
            .O(N__27007),
            .I(N__26997));
    InMux I__3731 (
            .O(N__27006),
            .I(N__26994));
    LocalMux I__3730 (
            .O(N__27003),
            .I(N__26991));
    Span4Mux_v I__3729 (
            .O(N__27000),
            .I(N__26988));
    LocalMux I__3728 (
            .O(N__26997),
            .I(N__26983));
    LocalMux I__3727 (
            .O(N__26994),
            .I(N__26983));
    Odrv4 I__3726 (
            .O(N__26991),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__3725 (
            .O(N__26988),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv12 I__3724 (
            .O(N__26983),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__3723 (
            .O(N__26976),
            .I(N__26973));
    LocalMux I__3722 (
            .O(N__26973),
            .I(N__26969));
    InMux I__3721 (
            .O(N__26972),
            .I(N__26966));
    Span4Mux_v I__3720 (
            .O(N__26969),
            .I(N__26959));
    LocalMux I__3719 (
            .O(N__26966),
            .I(N__26959));
    InMux I__3718 (
            .O(N__26965),
            .I(N__26954));
    InMux I__3717 (
            .O(N__26964),
            .I(N__26954));
    Span4Mux_v I__3716 (
            .O(N__26959),
            .I(N__26951));
    LocalMux I__3715 (
            .O(N__26954),
            .I(N__26948));
    Odrv4 I__3714 (
            .O(N__26951),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv12 I__3713 (
            .O(N__26948),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__3712 (
            .O(N__26943),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__3711 (
            .O(N__26940),
            .I(N__26936));
    InMux I__3710 (
            .O(N__26939),
            .I(N__26932));
    InMux I__3709 (
            .O(N__26936),
            .I(N__26929));
    InMux I__3708 (
            .O(N__26935),
            .I(N__26926));
    LocalMux I__3707 (
            .O(N__26932),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    LocalMux I__3706 (
            .O(N__26929),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    LocalMux I__3705 (
            .O(N__26926),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__3704 (
            .O(N__26919),
            .I(N__26913));
    InMux I__3703 (
            .O(N__26918),
            .I(N__26910));
    InMux I__3702 (
            .O(N__26917),
            .I(N__26907));
    InMux I__3701 (
            .O(N__26916),
            .I(N__26904));
    LocalMux I__3700 (
            .O(N__26913),
            .I(N__26901));
    LocalMux I__3699 (
            .O(N__26910),
            .I(N__26894));
    LocalMux I__3698 (
            .O(N__26907),
            .I(N__26894));
    LocalMux I__3697 (
            .O(N__26904),
            .I(N__26894));
    Odrv4 I__3696 (
            .O(N__26901),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv12 I__3695 (
            .O(N__26894),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__3694 (
            .O(N__26889),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__3693 (
            .O(N__26886),
            .I(N__26882));
    InMux I__3692 (
            .O(N__26885),
            .I(N__26878));
    InMux I__3691 (
            .O(N__26882),
            .I(N__26875));
    InMux I__3690 (
            .O(N__26881),
            .I(N__26872));
    LocalMux I__3689 (
            .O(N__26878),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    LocalMux I__3688 (
            .O(N__26875),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    LocalMux I__3687 (
            .O(N__26872),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    CascadeMux I__3686 (
            .O(N__26865),
            .I(N__26862));
    InMux I__3685 (
            .O(N__26862),
            .I(N__26858));
    InMux I__3684 (
            .O(N__26861),
            .I(N__26853));
    LocalMux I__3683 (
            .O(N__26858),
            .I(N__26850));
    InMux I__3682 (
            .O(N__26857),
            .I(N__26847));
    InMux I__3681 (
            .O(N__26856),
            .I(N__26844));
    LocalMux I__3680 (
            .O(N__26853),
            .I(N__26841));
    Sp12to4 I__3679 (
            .O(N__26850),
            .I(N__26834));
    LocalMux I__3678 (
            .O(N__26847),
            .I(N__26834));
    LocalMux I__3677 (
            .O(N__26844),
            .I(N__26834));
    Odrv4 I__3676 (
            .O(N__26841),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv12 I__3675 (
            .O(N__26834),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__3674 (
            .O(N__26829),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__3673 (
            .O(N__26826),
            .I(N__26822));
    InMux I__3672 (
            .O(N__26825),
            .I(N__26818));
    InMux I__3671 (
            .O(N__26822),
            .I(N__26815));
    InMux I__3670 (
            .O(N__26821),
            .I(N__26812));
    LocalMux I__3669 (
            .O(N__26818),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    LocalMux I__3668 (
            .O(N__26815),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    LocalMux I__3667 (
            .O(N__26812),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    CascadeMux I__3666 (
            .O(N__26805),
            .I(N__26800));
    InMux I__3665 (
            .O(N__26804),
            .I(N__26796));
    CascadeMux I__3664 (
            .O(N__26803),
            .I(N__26793));
    InMux I__3663 (
            .O(N__26800),
            .I(N__26788));
    InMux I__3662 (
            .O(N__26799),
            .I(N__26788));
    LocalMux I__3661 (
            .O(N__26796),
            .I(N__26785));
    InMux I__3660 (
            .O(N__26793),
            .I(N__26782));
    LocalMux I__3659 (
            .O(N__26788),
            .I(N__26779));
    Span4Mux_v I__3658 (
            .O(N__26785),
            .I(N__26776));
    LocalMux I__3657 (
            .O(N__26782),
            .I(N__26771));
    Span4Mux_v I__3656 (
            .O(N__26779),
            .I(N__26771));
    Span4Mux_v I__3655 (
            .O(N__26776),
            .I(N__26768));
    Odrv4 I__3654 (
            .O(N__26771),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__3653 (
            .O(N__26768),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__3652 (
            .O(N__26763),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__3651 (
            .O(N__26760),
            .I(N__26756));
    InMux I__3650 (
            .O(N__26759),
            .I(N__26752));
    InMux I__3649 (
            .O(N__26756),
            .I(N__26749));
    InMux I__3648 (
            .O(N__26755),
            .I(N__26746));
    LocalMux I__3647 (
            .O(N__26752),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    LocalMux I__3646 (
            .O(N__26749),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    LocalMux I__3645 (
            .O(N__26746),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    CascadeMux I__3644 (
            .O(N__26739),
            .I(N__26736));
    InMux I__3643 (
            .O(N__26736),
            .I(N__26731));
    InMux I__3642 (
            .O(N__26735),
            .I(N__26727));
    InMux I__3641 (
            .O(N__26734),
            .I(N__26724));
    LocalMux I__3640 (
            .O(N__26731),
            .I(N__26721));
    InMux I__3639 (
            .O(N__26730),
            .I(N__26718));
    LocalMux I__3638 (
            .O(N__26727),
            .I(N__26713));
    LocalMux I__3637 (
            .O(N__26724),
            .I(N__26713));
    Span4Mux_v I__3636 (
            .O(N__26721),
            .I(N__26706));
    LocalMux I__3635 (
            .O(N__26718),
            .I(N__26706));
    Span4Mux_h I__3634 (
            .O(N__26713),
            .I(N__26706));
    Span4Mux_v I__3633 (
            .O(N__26706),
            .I(N__26703));
    Odrv4 I__3632 (
            .O(N__26703),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__3631 (
            .O(N__26700),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__3630 (
            .O(N__26697),
            .I(N__26693));
    InMux I__3629 (
            .O(N__26696),
            .I(N__26689));
    InMux I__3628 (
            .O(N__26693),
            .I(N__26686));
    InMux I__3627 (
            .O(N__26692),
            .I(N__26683));
    LocalMux I__3626 (
            .O(N__26689),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    LocalMux I__3625 (
            .O(N__26686),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    LocalMux I__3624 (
            .O(N__26683),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__3623 (
            .O(N__26676),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__3622 (
            .O(N__26673),
            .I(N__26670));
    InMux I__3621 (
            .O(N__26670),
            .I(N__26667));
    LocalMux I__3620 (
            .O(N__26667),
            .I(N__26664));
    Odrv12 I__3619 (
            .O(N__26664),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__3618 (
            .O(N__26661),
            .I(N__26658));
    LocalMux I__3617 (
            .O(N__26658),
            .I(N__26655));
    Odrv4 I__3616 (
            .O(N__26655),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__3615 (
            .O(N__26652),
            .I(N__26649));
    LocalMux I__3614 (
            .O(N__26649),
            .I(N__26646));
    Span4Mux_v I__3613 (
            .O(N__26646),
            .I(N__26643));
    Odrv4 I__3612 (
            .O(N__26643),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    CascadeMux I__3611 (
            .O(N__26640),
            .I(N__26637));
    InMux I__3610 (
            .O(N__26637),
            .I(N__26634));
    LocalMux I__3609 (
            .O(N__26634),
            .I(N__26631));
    Span4Mux_h I__3608 (
            .O(N__26631),
            .I(N__26628));
    Odrv4 I__3607 (
            .O(N__26628),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    CascadeMux I__3606 (
            .O(N__26625),
            .I(N__26622));
    InMux I__3605 (
            .O(N__26622),
            .I(N__26619));
    LocalMux I__3604 (
            .O(N__26619),
            .I(N__26616));
    Span4Mux_v I__3603 (
            .O(N__26616),
            .I(N__26613));
    Odrv4 I__3602 (
            .O(N__26613),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__3601 (
            .O(N__26610),
            .I(N__26607));
    InMux I__3600 (
            .O(N__26607),
            .I(N__26604));
    LocalMux I__3599 (
            .O(N__26604),
            .I(N__26601));
    Odrv4 I__3598 (
            .O(N__26601),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    CascadeMux I__3597 (
            .O(N__26598),
            .I(N__26595));
    InMux I__3596 (
            .O(N__26595),
            .I(N__26592));
    LocalMux I__3595 (
            .O(N__26592),
            .I(N__26589));
    Span4Mux_h I__3594 (
            .O(N__26589),
            .I(N__26586));
    Odrv4 I__3593 (
            .O(N__26586),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__3592 (
            .O(N__26583),
            .I(N__26580));
    InMux I__3591 (
            .O(N__26580),
            .I(N__26577));
    LocalMux I__3590 (
            .O(N__26577),
            .I(N__26574));
    Span4Mux_h I__3589 (
            .O(N__26574),
            .I(N__26571));
    Odrv4 I__3588 (
            .O(N__26571),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__3587 (
            .O(N__26568),
            .I(N__26565));
    InMux I__3586 (
            .O(N__26565),
            .I(N__26562));
    LocalMux I__3585 (
            .O(N__26562),
            .I(N__26559));
    Odrv4 I__3584 (
            .O(N__26559),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__3583 (
            .O(N__26556),
            .I(N__26553));
    LocalMux I__3582 (
            .O(N__26553),
            .I(N__26550));
    Span4Mux_h I__3581 (
            .O(N__26550),
            .I(N__26547));
    Odrv4 I__3580 (
            .O(N__26547),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__3579 (
            .O(N__26544),
            .I(N__26541));
    LocalMux I__3578 (
            .O(N__26541),
            .I(N__26538));
    Span4Mux_v I__3577 (
            .O(N__26538),
            .I(N__26535));
    Odrv4 I__3576 (
            .O(N__26535),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    CascadeMux I__3575 (
            .O(N__26532),
            .I(N__26529));
    InMux I__3574 (
            .O(N__26529),
            .I(N__26526));
    LocalMux I__3573 (
            .O(N__26526),
            .I(N__26523));
    Odrv12 I__3572 (
            .O(N__26523),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__3571 (
            .O(N__26520),
            .I(N__26517));
    InMux I__3570 (
            .O(N__26517),
            .I(N__26514));
    LocalMux I__3569 (
            .O(N__26514),
            .I(N__26511));
    Span4Mux_h I__3568 (
            .O(N__26511),
            .I(N__26508));
    Span4Mux_h I__3567 (
            .O(N__26508),
            .I(N__26505));
    Odrv4 I__3566 (
            .O(N__26505),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__3565 (
            .O(N__26502),
            .I(N__26499));
    InMux I__3564 (
            .O(N__26499),
            .I(N__26496));
    LocalMux I__3563 (
            .O(N__26496),
            .I(N__26493));
    Odrv4 I__3562 (
            .O(N__26493),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    CascadeMux I__3561 (
            .O(N__26490),
            .I(N__26487));
    InMux I__3560 (
            .O(N__26487),
            .I(N__26484));
    LocalMux I__3559 (
            .O(N__26484),
            .I(N__26481));
    Odrv4 I__3558 (
            .O(N__26481),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__3557 (
            .O(N__26478),
            .I(N__26475));
    InMux I__3556 (
            .O(N__26475),
            .I(N__26472));
    LocalMux I__3555 (
            .O(N__26472),
            .I(N__26469));
    Span4Mux_h I__3554 (
            .O(N__26469),
            .I(N__26466));
    Odrv4 I__3553 (
            .O(N__26466),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    CascadeMux I__3552 (
            .O(N__26463),
            .I(N__26460));
    InMux I__3551 (
            .O(N__26460),
            .I(N__26457));
    LocalMux I__3550 (
            .O(N__26457),
            .I(N__26454));
    Span4Mux_h I__3549 (
            .O(N__26454),
            .I(N__26451));
    Odrv4 I__3548 (
            .O(N__26451),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    CascadeMux I__3547 (
            .O(N__26448),
            .I(N__26445));
    InMux I__3546 (
            .O(N__26445),
            .I(N__26442));
    LocalMux I__3545 (
            .O(N__26442),
            .I(N__26439));
    Odrv4 I__3544 (
            .O(N__26439),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__3543 (
            .O(N__26436),
            .I(N__26433));
    InMux I__3542 (
            .O(N__26433),
            .I(N__26430));
    LocalMux I__3541 (
            .O(N__26430),
            .I(N__26427));
    Odrv4 I__3540 (
            .O(N__26427),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__3539 (
            .O(N__26424),
            .I(N__26421));
    InMux I__3538 (
            .O(N__26421),
            .I(N__26418));
    LocalMux I__3537 (
            .O(N__26418),
            .I(N__26415));
    Span4Mux_v I__3536 (
            .O(N__26415),
            .I(N__26412));
    Odrv4 I__3535 (
            .O(N__26412),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__3534 (
            .O(N__26409),
            .I(N__26406));
    LocalMux I__3533 (
            .O(N__26406),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__3532 (
            .O(N__26403),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__3531 (
            .O(N__26400),
            .I(N__26396));
    CascadeMux I__3530 (
            .O(N__26399),
            .I(N__26393));
    LocalMux I__3529 (
            .O(N__26396),
            .I(N__26390));
    InMux I__3528 (
            .O(N__26393),
            .I(N__26387));
    Span4Mux_v I__3527 (
            .O(N__26390),
            .I(N__26382));
    LocalMux I__3526 (
            .O(N__26387),
            .I(N__26382));
    Span4Mux_v I__3525 (
            .O(N__26382),
            .I(N__26379));
    Span4Mux_v I__3524 (
            .O(N__26379),
            .I(N__26376));
    Odrv4 I__3523 (
            .O(N__26376),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__3522 (
            .O(N__26373),
            .I(N__26370));
    LocalMux I__3521 (
            .O(N__26370),
            .I(N__26367));
    Span4Mux_h I__3520 (
            .O(N__26367),
            .I(N__26364));
    Span4Mux_v I__3519 (
            .O(N__26364),
            .I(N__26361));
    Odrv4 I__3518 (
            .O(N__26361),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    CascadeMux I__3517 (
            .O(N__26358),
            .I(N__26355));
    InMux I__3516 (
            .O(N__26355),
            .I(N__26352));
    LocalMux I__3515 (
            .O(N__26352),
            .I(N__26349));
    Span4Mux_h I__3514 (
            .O(N__26349),
            .I(N__26346));
    Span4Mux_h I__3513 (
            .O(N__26346),
            .I(N__26343));
    Odrv4 I__3512 (
            .O(N__26343),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    CascadeMux I__3511 (
            .O(N__26340),
            .I(N__26337));
    InMux I__3510 (
            .O(N__26337),
            .I(N__26334));
    LocalMux I__3509 (
            .O(N__26334),
            .I(N__26331));
    Span4Mux_v I__3508 (
            .O(N__26331),
            .I(N__26328));
    Odrv4 I__3507 (
            .O(N__26328),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__3506 (
            .O(N__26325),
            .I(N__26322));
    LocalMux I__3505 (
            .O(N__26322),
            .I(N__26319));
    Odrv4 I__3504 (
            .O(N__26319),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    CascadeMux I__3503 (
            .O(N__26316),
            .I(N__26313));
    InMux I__3502 (
            .O(N__26313),
            .I(N__26310));
    LocalMux I__3501 (
            .O(N__26310),
            .I(N__26307));
    Span4Mux_h I__3500 (
            .O(N__26307),
            .I(N__26304));
    Odrv4 I__3499 (
            .O(N__26304),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__3498 (
            .O(N__26301),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_28 ));
    InMux I__3497 (
            .O(N__26298),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_29 ));
    InMux I__3496 (
            .O(N__26295),
            .I(N__26255));
    InMux I__3495 (
            .O(N__26294),
            .I(N__26255));
    InMux I__3494 (
            .O(N__26293),
            .I(N__26255));
    InMux I__3493 (
            .O(N__26292),
            .I(N__26255));
    InMux I__3492 (
            .O(N__26291),
            .I(N__26246));
    InMux I__3491 (
            .O(N__26290),
            .I(N__26246));
    InMux I__3490 (
            .O(N__26289),
            .I(N__26246));
    InMux I__3489 (
            .O(N__26288),
            .I(N__26246));
    InMux I__3488 (
            .O(N__26287),
            .I(N__26237));
    InMux I__3487 (
            .O(N__26286),
            .I(N__26237));
    InMux I__3486 (
            .O(N__26285),
            .I(N__26237));
    InMux I__3485 (
            .O(N__26284),
            .I(N__26237));
    InMux I__3484 (
            .O(N__26283),
            .I(N__26228));
    InMux I__3483 (
            .O(N__26282),
            .I(N__26228));
    InMux I__3482 (
            .O(N__26281),
            .I(N__26228));
    InMux I__3481 (
            .O(N__26280),
            .I(N__26228));
    InMux I__3480 (
            .O(N__26279),
            .I(N__26219));
    InMux I__3479 (
            .O(N__26278),
            .I(N__26219));
    InMux I__3478 (
            .O(N__26277),
            .I(N__26219));
    InMux I__3477 (
            .O(N__26276),
            .I(N__26219));
    InMux I__3476 (
            .O(N__26275),
            .I(N__26210));
    InMux I__3475 (
            .O(N__26274),
            .I(N__26210));
    InMux I__3474 (
            .O(N__26273),
            .I(N__26210));
    InMux I__3473 (
            .O(N__26272),
            .I(N__26210));
    InMux I__3472 (
            .O(N__26271),
            .I(N__26201));
    InMux I__3471 (
            .O(N__26270),
            .I(N__26201));
    InMux I__3470 (
            .O(N__26269),
            .I(N__26201));
    InMux I__3469 (
            .O(N__26268),
            .I(N__26201));
    InMux I__3468 (
            .O(N__26267),
            .I(N__26192));
    InMux I__3467 (
            .O(N__26266),
            .I(N__26192));
    InMux I__3466 (
            .O(N__26265),
            .I(N__26192));
    InMux I__3465 (
            .O(N__26264),
            .I(N__26192));
    LocalMux I__3464 (
            .O(N__26255),
            .I(N__26183));
    LocalMux I__3463 (
            .O(N__26246),
            .I(N__26183));
    LocalMux I__3462 (
            .O(N__26237),
            .I(N__26183));
    LocalMux I__3461 (
            .O(N__26228),
            .I(N__26183));
    LocalMux I__3460 (
            .O(N__26219),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__3459 (
            .O(N__26210),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__3458 (
            .O(N__26201),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__3457 (
            .O(N__26192),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    Odrv4 I__3456 (
            .O(N__26183),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    InMux I__3455 (
            .O(N__26172),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_30 ));
    CEMux I__3454 (
            .O(N__26169),
            .I(N__26157));
    CEMux I__3453 (
            .O(N__26168),
            .I(N__26157));
    CEMux I__3452 (
            .O(N__26167),
            .I(N__26157));
    CEMux I__3451 (
            .O(N__26166),
            .I(N__26157));
    GlobalMux I__3450 (
            .O(N__26157),
            .I(N__26154));
    gio2CtrlBuf I__3449 (
            .O(N__26154),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_g ));
    InMux I__3448 (
            .O(N__26151),
            .I(N__26147));
    InMux I__3447 (
            .O(N__26150),
            .I(N__26144));
    LocalMux I__3446 (
            .O(N__26147),
            .I(N__26141));
    LocalMux I__3445 (
            .O(N__26144),
            .I(N__26138));
    Span4Mux_v I__3444 (
            .O(N__26141),
            .I(N__26135));
    Span4Mux_v I__3443 (
            .O(N__26138),
            .I(N__26132));
    Span4Mux_h I__3442 (
            .O(N__26135),
            .I(N__26129));
    Span4Mux_h I__3441 (
            .O(N__26132),
            .I(N__26126));
    Odrv4 I__3440 (
            .O(N__26129),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__3439 (
            .O(N__26126),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__3438 (
            .O(N__26121),
            .I(N__26118));
    LocalMux I__3437 (
            .O(N__26118),
            .I(N__26114));
    InMux I__3436 (
            .O(N__26117),
            .I(N__26111));
    Sp12to4 I__3435 (
            .O(N__26114),
            .I(N__26106));
    LocalMux I__3434 (
            .O(N__26111),
            .I(N__26106));
    Odrv12 I__3433 (
            .O(N__26106),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__3432 (
            .O(N__26103),
            .I(N__26099));
    InMux I__3431 (
            .O(N__26102),
            .I(N__26096));
    LocalMux I__3430 (
            .O(N__26099),
            .I(N__26093));
    LocalMux I__3429 (
            .O(N__26096),
            .I(N__26090));
    Span12Mux_s5_h I__3428 (
            .O(N__26093),
            .I(N__26087));
    Odrv12 I__3427 (
            .O(N__26090),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    Odrv12 I__3426 (
            .O(N__26087),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__3425 (
            .O(N__26082),
            .I(N__26078));
    InMux I__3424 (
            .O(N__26081),
            .I(N__26075));
    LocalMux I__3423 (
            .O(N__26078),
            .I(N__26072));
    LocalMux I__3422 (
            .O(N__26075),
            .I(N__26069));
    Span4Mux_s3_h I__3421 (
            .O(N__26072),
            .I(N__26066));
    Odrv12 I__3420 (
            .O(N__26069),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv4 I__3419 (
            .O(N__26066),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__3418 (
            .O(N__26061),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_19 ));
    InMux I__3417 (
            .O(N__26058),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_20 ));
    InMux I__3416 (
            .O(N__26055),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_21 ));
    InMux I__3415 (
            .O(N__26052),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_22 ));
    InMux I__3414 (
            .O(N__26049),
            .I(bfn_10_10_0_));
    InMux I__3413 (
            .O(N__26046),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_24 ));
    InMux I__3412 (
            .O(N__26043),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_25 ));
    InMux I__3411 (
            .O(N__26040),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_26 ));
    InMux I__3410 (
            .O(N__26037),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_27 ));
    InMux I__3409 (
            .O(N__26034),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_10 ));
    InMux I__3408 (
            .O(N__26031),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_11 ));
    InMux I__3407 (
            .O(N__26028),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_12 ));
    InMux I__3406 (
            .O(N__26025),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_13 ));
    InMux I__3405 (
            .O(N__26022),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_14 ));
    InMux I__3404 (
            .O(N__26019),
            .I(bfn_10_9_0_));
    InMux I__3403 (
            .O(N__26016),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_16 ));
    InMux I__3402 (
            .O(N__26013),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_17 ));
    InMux I__3401 (
            .O(N__26010),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_18 ));
    InMux I__3400 (
            .O(N__26007),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_1 ));
    InMux I__3399 (
            .O(N__26004),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_2 ));
    InMux I__3398 (
            .O(N__26001),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_3 ));
    InMux I__3397 (
            .O(N__25998),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_4 ));
    InMux I__3396 (
            .O(N__25995),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_5 ));
    InMux I__3395 (
            .O(N__25992),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_6 ));
    InMux I__3394 (
            .O(N__25989),
            .I(bfn_10_8_0_));
    InMux I__3393 (
            .O(N__25986),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_8 ));
    InMux I__3392 (
            .O(N__25983),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_9 ));
    InMux I__3391 (
            .O(N__25980),
            .I(N__25977));
    LocalMux I__3390 (
            .O(N__25977),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__3389 (
            .O(N__25974),
            .I(N__25948));
    InMux I__3388 (
            .O(N__25973),
            .I(N__25948));
    InMux I__3387 (
            .O(N__25972),
            .I(N__25935));
    InMux I__3386 (
            .O(N__25971),
            .I(N__25935));
    InMux I__3385 (
            .O(N__25970),
            .I(N__25935));
    InMux I__3384 (
            .O(N__25969),
            .I(N__25935));
    InMux I__3383 (
            .O(N__25968),
            .I(N__25922));
    InMux I__3382 (
            .O(N__25967),
            .I(N__25922));
    InMux I__3381 (
            .O(N__25966),
            .I(N__25922));
    InMux I__3380 (
            .O(N__25965),
            .I(N__25922));
    InMux I__3379 (
            .O(N__25964),
            .I(N__25913));
    InMux I__3378 (
            .O(N__25963),
            .I(N__25913));
    InMux I__3377 (
            .O(N__25962),
            .I(N__25913));
    InMux I__3376 (
            .O(N__25961),
            .I(N__25913));
    InMux I__3375 (
            .O(N__25960),
            .I(N__25904));
    InMux I__3374 (
            .O(N__25959),
            .I(N__25904));
    InMux I__3373 (
            .O(N__25958),
            .I(N__25904));
    InMux I__3372 (
            .O(N__25957),
            .I(N__25904));
    InMux I__3371 (
            .O(N__25956),
            .I(N__25895));
    InMux I__3370 (
            .O(N__25955),
            .I(N__25895));
    InMux I__3369 (
            .O(N__25954),
            .I(N__25895));
    InMux I__3368 (
            .O(N__25953),
            .I(N__25895));
    LocalMux I__3367 (
            .O(N__25948),
            .I(N__25892));
    InMux I__3366 (
            .O(N__25947),
            .I(N__25883));
    InMux I__3365 (
            .O(N__25946),
            .I(N__25883));
    InMux I__3364 (
            .O(N__25945),
            .I(N__25883));
    InMux I__3363 (
            .O(N__25944),
            .I(N__25883));
    LocalMux I__3362 (
            .O(N__25935),
            .I(N__25880));
    InMux I__3361 (
            .O(N__25934),
            .I(N__25871));
    InMux I__3360 (
            .O(N__25933),
            .I(N__25871));
    InMux I__3359 (
            .O(N__25932),
            .I(N__25871));
    InMux I__3358 (
            .O(N__25931),
            .I(N__25871));
    LocalMux I__3357 (
            .O(N__25922),
            .I(N__25862));
    LocalMux I__3356 (
            .O(N__25913),
            .I(N__25862));
    LocalMux I__3355 (
            .O(N__25904),
            .I(N__25862));
    LocalMux I__3354 (
            .O(N__25895),
            .I(N__25862));
    Span4Mux_v I__3353 (
            .O(N__25892),
            .I(N__25857));
    LocalMux I__3352 (
            .O(N__25883),
            .I(N__25857));
    Span4Mux_v I__3351 (
            .O(N__25880),
            .I(N__25848));
    LocalMux I__3350 (
            .O(N__25871),
            .I(N__25848));
    Span4Mux_v I__3349 (
            .O(N__25862),
            .I(N__25848));
    Span4Mux_h I__3348 (
            .O(N__25857),
            .I(N__25848));
    Odrv4 I__3347 (
            .O(N__25848),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__3346 (
            .O(N__25845),
            .I(N__25842));
    LocalMux I__3345 (
            .O(N__25842),
            .I(N__25837));
    InMux I__3344 (
            .O(N__25841),
            .I(N__25832));
    InMux I__3343 (
            .O(N__25840),
            .I(N__25832));
    Span12Mux_s11_v I__3342 (
            .O(N__25837),
            .I(N__25828));
    LocalMux I__3341 (
            .O(N__25832),
            .I(N__25825));
    InMux I__3340 (
            .O(N__25831),
            .I(N__25822));
    Span12Mux_v I__3339 (
            .O(N__25828),
            .I(N__25819));
    Odrv4 I__3338 (
            .O(N__25825),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__3337 (
            .O(N__25822),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__3336 (
            .O(N__25819),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__3335 (
            .O(N__25812),
            .I(N__25809));
    LocalMux I__3334 (
            .O(N__25809),
            .I(N__25806));
    Odrv12 I__3333 (
            .O(N__25806),
            .I(s3_phy_c));
    CascadeMux I__3332 (
            .O(N__25803),
            .I(N__25798));
    InMux I__3331 (
            .O(N__25802),
            .I(N__25790));
    InMux I__3330 (
            .O(N__25801),
            .I(N__25790));
    InMux I__3329 (
            .O(N__25798),
            .I(N__25790));
    InMux I__3328 (
            .O(N__25797),
            .I(N__25787));
    LocalMux I__3327 (
            .O(N__25790),
            .I(N__25782));
    LocalMux I__3326 (
            .O(N__25787),
            .I(N__25782));
    Odrv4 I__3325 (
            .O(N__25782),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__3324 (
            .O(N__25779),
            .I(N__25776));
    LocalMux I__3323 (
            .O(N__25776),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__3322 (
            .O(N__25773),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_0 ));
    InMux I__3321 (
            .O(N__25770),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__3320 (
            .O(N__25767),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__3319 (
            .O(N__25764),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__3318 (
            .O(N__25761),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__3317 (
            .O(N__25758),
            .I(bfn_9_22_0_));
    InMux I__3316 (
            .O(N__25755),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__3315 (
            .O(N__25752),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__3314 (
            .O(N__25749),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__3313 (
            .O(N__25746),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__3312 (
            .O(N__25743),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__3311 (
            .O(N__25740),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__3310 (
            .O(N__25737),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__3309 (
            .O(N__25734),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__3308 (
            .O(N__25731),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__3307 (
            .O(N__25728),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__3306 (
            .O(N__25725),
            .I(bfn_9_21_0_));
    InMux I__3305 (
            .O(N__25722),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__3304 (
            .O(N__25719),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__3303 (
            .O(N__25716),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__3302 (
            .O(N__25713),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__3301 (
            .O(N__25710),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__3300 (
            .O(N__25707),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    InMux I__3299 (
            .O(N__25704),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__3298 (
            .O(N__25701),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__3297 (
            .O(N__25698),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__3296 (
            .O(N__25695),
            .I(bfn_9_20_0_));
    InMux I__3295 (
            .O(N__25692),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__3294 (
            .O(N__25689),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__3293 (
            .O(N__25686),
            .I(N__25683));
    LocalMux I__3292 (
            .O(N__25683),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__3291 (
            .O(N__25680),
            .I(N__25677));
    InMux I__3290 (
            .O(N__25677),
            .I(N__25674));
    LocalMux I__3289 (
            .O(N__25674),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    CascadeMux I__3288 (
            .O(N__25671),
            .I(N__25668));
    InMux I__3287 (
            .O(N__25668),
            .I(N__25665));
    LocalMux I__3286 (
            .O(N__25665),
            .I(N__25662));
    Span4Mux_v I__3285 (
            .O(N__25662),
            .I(N__25658));
    InMux I__3284 (
            .O(N__25661),
            .I(N__25653));
    Span4Mux_v I__3283 (
            .O(N__25658),
            .I(N__25650));
    InMux I__3282 (
            .O(N__25657),
            .I(N__25647));
    InMux I__3281 (
            .O(N__25656),
            .I(N__25644));
    LocalMux I__3280 (
            .O(N__25653),
            .I(N__25641));
    Odrv4 I__3279 (
            .O(N__25650),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__3278 (
            .O(N__25647),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__3277 (
            .O(N__25644),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv12 I__3276 (
            .O(N__25641),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__3275 (
            .O(N__25632),
            .I(N__25629));
    InMux I__3274 (
            .O(N__25629),
            .I(N__25626));
    LocalMux I__3273 (
            .O(N__25626),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__3272 (
            .O(N__25623),
            .I(N__25620));
    LocalMux I__3271 (
            .O(N__25620),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    CascadeMux I__3270 (
            .O(N__25617),
            .I(N__25614));
    InMux I__3269 (
            .O(N__25614),
            .I(N__25611));
    LocalMux I__3268 (
            .O(N__25611),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__3267 (
            .O(N__25608),
            .I(N__25605));
    LocalMux I__3266 (
            .O(N__25605),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__3265 (
            .O(N__25602),
            .I(N__25599));
    InMux I__3264 (
            .O(N__25599),
            .I(N__25596));
    LocalMux I__3263 (
            .O(N__25596),
            .I(N__25593));
    Odrv4 I__3262 (
            .O(N__25593),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__3261 (
            .O(N__25590),
            .I(bfn_9_19_0_));
    InMux I__3260 (
            .O(N__25587),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__3259 (
            .O(N__25584),
            .I(N__25581));
    InMux I__3258 (
            .O(N__25581),
            .I(N__25578));
    LocalMux I__3257 (
            .O(N__25578),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__3256 (
            .O(N__25575),
            .I(N__25572));
    LocalMux I__3255 (
            .O(N__25572),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__3254 (
            .O(N__25569),
            .I(N__25566));
    LocalMux I__3253 (
            .O(N__25566),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__3252 (
            .O(N__25563),
            .I(N__25560));
    LocalMux I__3251 (
            .O(N__25560),
            .I(N__25557));
    Span4Mux_h I__3250 (
            .O(N__25557),
            .I(N__25554));
    Odrv4 I__3249 (
            .O(N__25554),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__3248 (
            .O(N__25551),
            .I(N__25548));
    LocalMux I__3247 (
            .O(N__25548),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__3246 (
            .O(N__25545),
            .I(N__25542));
    InMux I__3245 (
            .O(N__25542),
            .I(N__25539));
    LocalMux I__3244 (
            .O(N__25539),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__3243 (
            .O(N__25536),
            .I(N__25533));
    InMux I__3242 (
            .O(N__25533),
            .I(N__25530));
    LocalMux I__3241 (
            .O(N__25530),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__3240 (
            .O(N__25527),
            .I(N__25524));
    InMux I__3239 (
            .O(N__25524),
            .I(N__25521));
    LocalMux I__3238 (
            .O(N__25521),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__3237 (
            .O(N__25518),
            .I(N__25515));
    InMux I__3236 (
            .O(N__25515),
            .I(N__25512));
    LocalMux I__3235 (
            .O(N__25512),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__3234 (
            .O(N__25509),
            .I(N__25506));
    LocalMux I__3233 (
            .O(N__25506),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__3232 (
            .O(N__25503),
            .I(N__25500));
    LocalMux I__3231 (
            .O(N__25500),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__3230 (
            .O(N__25497),
            .I(N__25494));
    LocalMux I__3229 (
            .O(N__25494),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__3228 (
            .O(N__25491),
            .I(N__25488));
    LocalMux I__3227 (
            .O(N__25488),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__3226 (
            .O(N__25485),
            .I(N__25482));
    LocalMux I__3225 (
            .O(N__25482),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__3224 (
            .O(N__25479),
            .I(N__25476));
    InMux I__3223 (
            .O(N__25476),
            .I(N__25473));
    LocalMux I__3222 (
            .O(N__25473),
            .I(N__25470));
    Span4Mux_v I__3221 (
            .O(N__25470),
            .I(N__25467));
    Odrv4 I__3220 (
            .O(N__25467),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    InMux I__3219 (
            .O(N__25464),
            .I(N__25461));
    LocalMux I__3218 (
            .O(N__25461),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__3217 (
            .O(N__25458),
            .I(N__25455));
    InMux I__3216 (
            .O(N__25455),
            .I(N__25452));
    LocalMux I__3215 (
            .O(N__25452),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__3214 (
            .O(N__25449),
            .I(N__25446));
    LocalMux I__3213 (
            .O(N__25446),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__3212 (
            .O(N__25443),
            .I(N__25440));
    InMux I__3211 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3210 (
            .O(N__25437),
            .I(N__25434));
    Odrv4 I__3209 (
            .O(N__25434),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__3208 (
            .O(N__25431),
            .I(N__25428));
    LocalMux I__3207 (
            .O(N__25428),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    CascadeMux I__3206 (
            .O(N__25425),
            .I(N__25422));
    InMux I__3205 (
            .O(N__25422),
            .I(N__25419));
    LocalMux I__3204 (
            .O(N__25419),
            .I(N__25416));
    Odrv4 I__3203 (
            .O(N__25416),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__3202 (
            .O(N__25413),
            .I(N__25410));
    InMux I__3201 (
            .O(N__25410),
            .I(N__25407));
    LocalMux I__3200 (
            .O(N__25407),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__3199 (
            .O(N__25404),
            .I(N__25401));
    LocalMux I__3198 (
            .O(N__25401),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__3197 (
            .O(N__25398),
            .I(N__25395));
    LocalMux I__3196 (
            .O(N__25395),
            .I(N__25392));
    Span4Mux_v I__3195 (
            .O(N__25392),
            .I(N__25389));
    Odrv4 I__3194 (
            .O(N__25389),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    CascadeMux I__3193 (
            .O(N__25386),
            .I(N__25383));
    InMux I__3192 (
            .O(N__25383),
            .I(N__25380));
    LocalMux I__3191 (
            .O(N__25380),
            .I(N__25377));
    Span4Mux_h I__3190 (
            .O(N__25377),
            .I(N__25374));
    Odrv4 I__3189 (
            .O(N__25374),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    CascadeMux I__3188 (
            .O(N__25371),
            .I(N__25368));
    InMux I__3187 (
            .O(N__25368),
            .I(N__25365));
    LocalMux I__3186 (
            .O(N__25365),
            .I(N__25362));
    Odrv4 I__3185 (
            .O(N__25362),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    CascadeMux I__3184 (
            .O(N__25359),
            .I(N__25356));
    InMux I__3183 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__3182 (
            .O(N__25353),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__3181 (
            .O(N__25350),
            .I(N__25347));
    LocalMux I__3180 (
            .O(N__25347),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    CascadeMux I__3179 (
            .O(N__25344),
            .I(N__25341));
    InMux I__3178 (
            .O(N__25341),
            .I(N__25338));
    LocalMux I__3177 (
            .O(N__25338),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__3176 (
            .O(N__25335),
            .I(N__25332));
    LocalMux I__3175 (
            .O(N__25332),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__3174 (
            .O(N__25329),
            .I(N__25326));
    LocalMux I__3173 (
            .O(N__25326),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    CascadeMux I__3172 (
            .O(N__25323),
            .I(N__25320));
    InMux I__3171 (
            .O(N__25320),
            .I(N__25317));
    LocalMux I__3170 (
            .O(N__25317),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__3169 (
            .O(N__25314),
            .I(N__25311));
    LocalMux I__3168 (
            .O(N__25311),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    CascadeMux I__3167 (
            .O(N__25308),
            .I(N__25305));
    InMux I__3166 (
            .O(N__25305),
            .I(N__25302));
    LocalMux I__3165 (
            .O(N__25302),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    CascadeMux I__3164 (
            .O(N__25299),
            .I(N__25296));
    InMux I__3163 (
            .O(N__25296),
            .I(N__25293));
    LocalMux I__3162 (
            .O(N__25293),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__3161 (
            .O(N__25290),
            .I(N__25287));
    LocalMux I__3160 (
            .O(N__25287),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__3159 (
            .O(N__25284),
            .I(N__25281));
    LocalMux I__3158 (
            .O(N__25281),
            .I(N__25277));
    CascadeMux I__3157 (
            .O(N__25280),
            .I(N__25274));
    Span12Mux_s8_v I__3156 (
            .O(N__25277),
            .I(N__25269));
    InMux I__3155 (
            .O(N__25274),
            .I(N__25266));
    InMux I__3154 (
            .O(N__25273),
            .I(N__25263));
    InMux I__3153 (
            .O(N__25272),
            .I(N__25260));
    Span12Mux_v I__3152 (
            .O(N__25269),
            .I(N__25257));
    LocalMux I__3151 (
            .O(N__25266),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3150 (
            .O(N__25263),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3149 (
            .O(N__25260),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__3148 (
            .O(N__25257),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__3147 (
            .O(N__25248),
            .I(N__25245));
    LocalMux I__3146 (
            .O(N__25245),
            .I(N__25242));
    Span4Mux_v I__3145 (
            .O(N__25242),
            .I(N__25237));
    InMux I__3144 (
            .O(N__25241),
            .I(N__25234));
    InMux I__3143 (
            .O(N__25240),
            .I(N__25231));
    Sp12to4 I__3142 (
            .O(N__25237),
            .I(N__25224));
    LocalMux I__3141 (
            .O(N__25234),
            .I(N__25224));
    LocalMux I__3140 (
            .O(N__25231),
            .I(N__25224));
    Span12Mux_h I__3139 (
            .O(N__25224),
            .I(N__25221));
    Odrv12 I__3138 (
            .O(N__25221),
            .I(il_min_comp2_c));
    CascadeMux I__3137 (
            .O(N__25218),
            .I(N__25213));
    InMux I__3136 (
            .O(N__25217),
            .I(N__25208));
    InMux I__3135 (
            .O(N__25216),
            .I(N__25208));
    InMux I__3134 (
            .O(N__25213),
            .I(N__25205));
    LocalMux I__3133 (
            .O(N__25208),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__3132 (
            .O(N__25205),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__3131 (
            .O(N__25200),
            .I(N__25197));
    InMux I__3130 (
            .O(N__25197),
            .I(N__25193));
    InMux I__3129 (
            .O(N__25196),
            .I(N__25190));
    LocalMux I__3128 (
            .O(N__25193),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__3127 (
            .O(N__25190),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    CascadeMux I__3126 (
            .O(N__25185),
            .I(N__25182));
    InMux I__3125 (
            .O(N__25182),
            .I(N__25179));
    LocalMux I__3124 (
            .O(N__25179),
            .I(\phase_controller_inst2.stoper_tr.un4_start_0 ));
    InMux I__3123 (
            .O(N__25176),
            .I(N__25173));
    LocalMux I__3122 (
            .O(N__25173),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__3121 (
            .O(N__25170),
            .I(N__25167));
    LocalMux I__3120 (
            .O(N__25167),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    CascadeMux I__3119 (
            .O(N__25164),
            .I(N__25161));
    InMux I__3118 (
            .O(N__25161),
            .I(N__25158));
    LocalMux I__3117 (
            .O(N__25158),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__3116 (
            .O(N__25155),
            .I(N__25152));
    LocalMux I__3115 (
            .O(N__25152),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__3114 (
            .O(N__25149),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__3113 (
            .O(N__25146),
            .I(N__25143));
    LocalMux I__3112 (
            .O(N__25143),
            .I(N__25140));
    Span4Mux_h I__3111 (
            .O(N__25140),
            .I(N__25137));
    Span4Mux_v I__3110 (
            .O(N__25137),
            .I(N__25134));
    Odrv4 I__3109 (
            .O(N__25134),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__3108 (
            .O(N__25131),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    CascadeMux I__3107 (
            .O(N__25128),
            .I(N__25125));
    InMux I__3106 (
            .O(N__25125),
            .I(N__25122));
    LocalMux I__3105 (
            .O(N__25122),
            .I(N__25119));
    Span4Mux_v I__3104 (
            .O(N__25119),
            .I(N__25116));
    Odrv4 I__3103 (
            .O(N__25116),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__3102 (
            .O(N__25113),
            .I(N__25110));
    LocalMux I__3101 (
            .O(N__25110),
            .I(N__25107));
    Span12Mux_v I__3100 (
            .O(N__25107),
            .I(N__25104));
    Odrv12 I__3099 (
            .O(N__25104),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__3098 (
            .O(N__25101),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__3097 (
            .O(N__25098),
            .I(N__25095));
    LocalMux I__3096 (
            .O(N__25095),
            .I(N__25092));
    Span4Mux_h I__3095 (
            .O(N__25092),
            .I(N__25089));
    Sp12to4 I__3094 (
            .O(N__25089),
            .I(N__25086));
    Odrv12 I__3093 (
            .O(N__25086),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__3092 (
            .O(N__25083),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__3091 (
            .O(N__25080),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__3090 (
            .O(N__25077),
            .I(N__25074));
    LocalMux I__3089 (
            .O(N__25074),
            .I(N__25071));
    Span12Mux_v I__3088 (
            .O(N__25071),
            .I(N__25068));
    Odrv12 I__3087 (
            .O(N__25068),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    CascadeMux I__3086 (
            .O(N__25065),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__3085 (
            .O(N__25062),
            .I(N__25059));
    LocalMux I__3084 (
            .O(N__25059),
            .I(N__25055));
    InMux I__3083 (
            .O(N__25058),
            .I(N__25052));
    Span12Mux_v I__3082 (
            .O(N__25055),
            .I(N__25047));
    LocalMux I__3081 (
            .O(N__25052),
            .I(N__25047));
    Odrv12 I__3080 (
            .O(N__25047),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    IoInMux I__3079 (
            .O(N__25044),
            .I(N__25041));
    LocalMux I__3078 (
            .O(N__25041),
            .I(N__25038));
    Odrv12 I__3077 (
            .O(N__25038),
            .I(s4_phy_c));
    InMux I__3076 (
            .O(N__25035),
            .I(N__25032));
    LocalMux I__3075 (
            .O(N__25032),
            .I(N__25029));
    Odrv4 I__3074 (
            .O(N__25029),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__3073 (
            .O(N__25026),
            .I(N__25023));
    LocalMux I__3072 (
            .O(N__25023),
            .I(N__25020));
    Span4Mux_h I__3071 (
            .O(N__25020),
            .I(N__25017));
    Odrv4 I__3070 (
            .O(N__25017),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__3069 (
            .O(N__25014),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    InMux I__3068 (
            .O(N__25011),
            .I(N__25008));
    LocalMux I__3067 (
            .O(N__25008),
            .I(N__25005));
    Sp12to4 I__3066 (
            .O(N__25005),
            .I(N__25002));
    Odrv12 I__3065 (
            .O(N__25002),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__3064 (
            .O(N__24999),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__3063 (
            .O(N__24996),
            .I(N__24993));
    LocalMux I__3062 (
            .O(N__24993),
            .I(N__24990));
    Span4Mux_h I__3061 (
            .O(N__24990),
            .I(N__24987));
    Sp12to4 I__3060 (
            .O(N__24987),
            .I(N__24984));
    Odrv12 I__3059 (
            .O(N__24984),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__3058 (
            .O(N__24981),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__3057 (
            .O(N__24978),
            .I(N__24975));
    LocalMux I__3056 (
            .O(N__24975),
            .I(N__24972));
    Span4Mux_v I__3055 (
            .O(N__24972),
            .I(N__24969));
    Odrv4 I__3054 (
            .O(N__24969),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__3053 (
            .O(N__24966),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__3052 (
            .O(N__24963),
            .I(N__24960));
    LocalMux I__3051 (
            .O(N__24960),
            .I(N__24957));
    Span4Mux_h I__3050 (
            .O(N__24957),
            .I(N__24954));
    Span4Mux_v I__3049 (
            .O(N__24954),
            .I(N__24951));
    Span4Mux_v I__3048 (
            .O(N__24951),
            .I(N__24948));
    Odrv4 I__3047 (
            .O(N__24948),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__3046 (
            .O(N__24945),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__3045 (
            .O(N__24942),
            .I(N__24939));
    LocalMux I__3044 (
            .O(N__24939),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__3043 (
            .O(N__24936),
            .I(N__24933));
    LocalMux I__3042 (
            .O(N__24933),
            .I(N__24930));
    Span4Mux_v I__3041 (
            .O(N__24930),
            .I(N__24927));
    Odrv4 I__3040 (
            .O(N__24927),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__3039 (
            .O(N__24924),
            .I(bfn_8_22_0_));
    InMux I__3038 (
            .O(N__24921),
            .I(N__24918));
    LocalMux I__3037 (
            .O(N__24918),
            .I(N__24915));
    Span4Mux_h I__3036 (
            .O(N__24915),
            .I(N__24912));
    Span4Mux_v I__3035 (
            .O(N__24912),
            .I(N__24909));
    Odrv4 I__3034 (
            .O(N__24909),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__3033 (
            .O(N__24906),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__3032 (
            .O(N__24903),
            .I(N__24900));
    LocalMux I__3031 (
            .O(N__24900),
            .I(N__24897));
    Span4Mux_h I__3030 (
            .O(N__24897),
            .I(N__24894));
    Span4Mux_v I__3029 (
            .O(N__24894),
            .I(N__24891));
    Span4Mux_h I__3028 (
            .O(N__24891),
            .I(N__24888));
    Odrv4 I__3027 (
            .O(N__24888),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__3026 (
            .O(N__24885),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__3025 (
            .O(N__24882),
            .I(N__24879));
    LocalMux I__3024 (
            .O(N__24879),
            .I(N__24876));
    Span4Mux_h I__3023 (
            .O(N__24876),
            .I(N__24873));
    Span4Mux_v I__3022 (
            .O(N__24873),
            .I(N__24870));
    Odrv4 I__3021 (
            .O(N__24870),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    CascadeMux I__3020 (
            .O(N__24867),
            .I(N__24864));
    InMux I__3019 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__3018 (
            .O(N__24861),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    InMux I__3017 (
            .O(N__24858),
            .I(N__24855));
    LocalMux I__3016 (
            .O(N__24855),
            .I(N__24852));
    Span4Mux_h I__3015 (
            .O(N__24852),
            .I(N__24849));
    Span4Mux_v I__3014 (
            .O(N__24849),
            .I(N__24846));
    Odrv4 I__3013 (
            .O(N__24846),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__3012 (
            .O(N__24843),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__3011 (
            .O(N__24840),
            .I(N__24837));
    LocalMux I__3010 (
            .O(N__24837),
            .I(N__24834));
    Sp12to4 I__3009 (
            .O(N__24834),
            .I(N__24831));
    Odrv12 I__3008 (
            .O(N__24831),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__3007 (
            .O(N__24828),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__3006 (
            .O(N__24825),
            .I(N__24822));
    LocalMux I__3005 (
            .O(N__24822),
            .I(N__24819));
    Span12Mux_s8_h I__3004 (
            .O(N__24819),
            .I(N__24816));
    Odrv12 I__3003 (
            .O(N__24816),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__3002 (
            .O(N__24813),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__3001 (
            .O(N__24810),
            .I(N__24807));
    LocalMux I__3000 (
            .O(N__24807),
            .I(N__24804));
    Span4Mux_v I__2999 (
            .O(N__24804),
            .I(N__24801));
    Span4Mux_v I__2998 (
            .O(N__24801),
            .I(N__24798));
    Odrv4 I__2997 (
            .O(N__24798),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__2996 (
            .O(N__24795),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__2995 (
            .O(N__24792),
            .I(N__24789));
    LocalMux I__2994 (
            .O(N__24789),
            .I(N__24786));
    Sp12to4 I__2993 (
            .O(N__24786),
            .I(N__24783));
    Span12Mux_v I__2992 (
            .O(N__24783),
            .I(N__24780));
    Odrv12 I__2991 (
            .O(N__24780),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__2990 (
            .O(N__24777),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__2989 (
            .O(N__24774),
            .I(N__24771));
    LocalMux I__2988 (
            .O(N__24771),
            .I(N__24768));
    Span12Mux_v I__2987 (
            .O(N__24768),
            .I(N__24765));
    Odrv12 I__2986 (
            .O(N__24765),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__2985 (
            .O(N__24762),
            .I(bfn_8_21_0_));
    InMux I__2984 (
            .O(N__24759),
            .I(N__24756));
    LocalMux I__2983 (
            .O(N__24756),
            .I(N__24753));
    Span4Mux_v I__2982 (
            .O(N__24753),
            .I(N__24750));
    Span4Mux_v I__2981 (
            .O(N__24750),
            .I(N__24747));
    Odrv4 I__2980 (
            .O(N__24747),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__2979 (
            .O(N__24744),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    CascadeMux I__2978 (
            .O(N__24741),
            .I(N__24738));
    InMux I__2977 (
            .O(N__24738),
            .I(N__24735));
    LocalMux I__2976 (
            .O(N__24735),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__2975 (
            .O(N__24732),
            .I(N__24729));
    LocalMux I__2974 (
            .O(N__24729),
            .I(N__24726));
    Span4Mux_v I__2973 (
            .O(N__24726),
            .I(N__24723));
    Odrv4 I__2972 (
            .O(N__24723),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__2971 (
            .O(N__24720),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__2970 (
            .O(N__24717),
            .I(N__24714));
    LocalMux I__2969 (
            .O(N__24714),
            .I(N__24711));
    Odrv4 I__2968 (
            .O(N__24711),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__2967 (
            .O(N__24708),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__2966 (
            .O(N__24705),
            .I(N__24702));
    LocalMux I__2965 (
            .O(N__24702),
            .I(N__24699));
    Odrv4 I__2964 (
            .O(N__24699),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__2963 (
            .O(N__24696),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__2962 (
            .O(N__24693),
            .I(N__24690));
    LocalMux I__2961 (
            .O(N__24690),
            .I(N__24687));
    Span12Mux_s8_h I__2960 (
            .O(N__24687),
            .I(N__24684));
    Odrv12 I__2959 (
            .O(N__24684),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__2958 (
            .O(N__24681),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    InMux I__2957 (
            .O(N__24678),
            .I(N__24675));
    LocalMux I__2956 (
            .O(N__24675),
            .I(N__24672));
    Odrv4 I__2955 (
            .O(N__24672),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__2954 (
            .O(N__24669),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__2953 (
            .O(N__24666),
            .I(N__24663));
    LocalMux I__2952 (
            .O(N__24663),
            .I(N__24660));
    Odrv4 I__2951 (
            .O(N__24660),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__2950 (
            .O(N__24657),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__2949 (
            .O(N__24654),
            .I(N__24651));
    LocalMux I__2948 (
            .O(N__24651),
            .I(N__24648));
    Span12Mux_v I__2947 (
            .O(N__24648),
            .I(N__24645));
    Odrv12 I__2946 (
            .O(N__24645),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__2945 (
            .O(N__24642),
            .I(bfn_8_20_0_));
    InMux I__2944 (
            .O(N__24639),
            .I(N__24636));
    LocalMux I__2943 (
            .O(N__24636),
            .I(N__24633));
    Span4Mux_h I__2942 (
            .O(N__24633),
            .I(N__24630));
    Span4Mux_v I__2941 (
            .O(N__24630),
            .I(N__24627));
    Odrv4 I__2940 (
            .O(N__24627),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__2939 (
            .O(N__24624),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__2938 (
            .O(N__24621),
            .I(N__24618));
    LocalMux I__2937 (
            .O(N__24618),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    InMux I__2936 (
            .O(N__24615),
            .I(N__24612));
    LocalMux I__2935 (
            .O(N__24612),
            .I(N__24609));
    Span4Mux_h I__2934 (
            .O(N__24609),
            .I(N__24606));
    Span4Mux_v I__2933 (
            .O(N__24606),
            .I(N__24603));
    Odrv4 I__2932 (
            .O(N__24603),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__2931 (
            .O(N__24600),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__2930 (
            .O(N__24597),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__2929 (
            .O(N__24594),
            .I(N__24589));
    InMux I__2928 (
            .O(N__24593),
            .I(N__24574));
    InMux I__2927 (
            .O(N__24592),
            .I(N__24574));
    InMux I__2926 (
            .O(N__24589),
            .I(N__24569));
    InMux I__2925 (
            .O(N__24588),
            .I(N__24569));
    CascadeMux I__2924 (
            .O(N__24587),
            .I(N__24566));
    InMux I__2923 (
            .O(N__24586),
            .I(N__24555));
    InMux I__2922 (
            .O(N__24585),
            .I(N__24544));
    InMux I__2921 (
            .O(N__24584),
            .I(N__24544));
    InMux I__2920 (
            .O(N__24583),
            .I(N__24544));
    InMux I__2919 (
            .O(N__24582),
            .I(N__24544));
    InMux I__2918 (
            .O(N__24581),
            .I(N__24544));
    CascadeMux I__2917 (
            .O(N__24580),
            .I(N__24541));
    CascadeMux I__2916 (
            .O(N__24579),
            .I(N__24537));
    LocalMux I__2915 (
            .O(N__24574),
            .I(N__24528));
    LocalMux I__2914 (
            .O(N__24569),
            .I(N__24528));
    InMux I__2913 (
            .O(N__24566),
            .I(N__24515));
    InMux I__2912 (
            .O(N__24565),
            .I(N__24515));
    InMux I__2911 (
            .O(N__24564),
            .I(N__24515));
    InMux I__2910 (
            .O(N__24563),
            .I(N__24515));
    InMux I__2909 (
            .O(N__24562),
            .I(N__24515));
    InMux I__2908 (
            .O(N__24561),
            .I(N__24515));
    InMux I__2907 (
            .O(N__24560),
            .I(N__24512));
    InMux I__2906 (
            .O(N__24559),
            .I(N__24509));
    InMux I__2905 (
            .O(N__24558),
            .I(N__24506));
    LocalMux I__2904 (
            .O(N__24555),
            .I(N__24501));
    LocalMux I__2903 (
            .O(N__24544),
            .I(N__24501));
    InMux I__2902 (
            .O(N__24541),
            .I(N__24496));
    InMux I__2901 (
            .O(N__24540),
            .I(N__24496));
    InMux I__2900 (
            .O(N__24537),
            .I(N__24493));
    InMux I__2899 (
            .O(N__24536),
            .I(N__24490));
    InMux I__2898 (
            .O(N__24535),
            .I(N__24483));
    InMux I__2897 (
            .O(N__24534),
            .I(N__24483));
    InMux I__2896 (
            .O(N__24533),
            .I(N__24483));
    Span4Mux_h I__2895 (
            .O(N__24528),
            .I(N__24476));
    LocalMux I__2894 (
            .O(N__24515),
            .I(N__24476));
    LocalMux I__2893 (
            .O(N__24512),
            .I(N__24476));
    LocalMux I__2892 (
            .O(N__24509),
            .I(N__24466));
    LocalMux I__2891 (
            .O(N__24506),
            .I(N__24466));
    Span4Mux_v I__2890 (
            .O(N__24501),
            .I(N__24466));
    LocalMux I__2889 (
            .O(N__24496),
            .I(N__24466));
    LocalMux I__2888 (
            .O(N__24493),
            .I(N__24459));
    LocalMux I__2887 (
            .O(N__24490),
            .I(N__24459));
    LocalMux I__2886 (
            .O(N__24483),
            .I(N__24459));
    Sp12to4 I__2885 (
            .O(N__24476),
            .I(N__24451));
    InMux I__2884 (
            .O(N__24475),
            .I(N__24448));
    Span4Mux_h I__2883 (
            .O(N__24466),
            .I(N__24443));
    Span4Mux_v I__2882 (
            .O(N__24459),
            .I(N__24443));
    InMux I__2881 (
            .O(N__24458),
            .I(N__24432));
    InMux I__2880 (
            .O(N__24457),
            .I(N__24432));
    InMux I__2879 (
            .O(N__24456),
            .I(N__24432));
    InMux I__2878 (
            .O(N__24455),
            .I(N__24432));
    InMux I__2877 (
            .O(N__24454),
            .I(N__24432));
    Span12Mux_v I__2876 (
            .O(N__24451),
            .I(N__24429));
    LocalMux I__2875 (
            .O(N__24448),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__2874 (
            .O(N__24443),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__2873 (
            .O(N__24432),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv12 I__2872 (
            .O(N__24429),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__2871 (
            .O(N__24420),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__2870 (
            .O(N__24417),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__2869 (
            .O(N__24414),
            .I(N__24411));
    LocalMux I__2868 (
            .O(N__24411),
            .I(N__24408));
    Odrv12 I__2867 (
            .O(N__24408),
            .I(\current_shift_inst.control_input_axb_28 ));
    CascadeMux I__2866 (
            .O(N__24405),
            .I(N__24402));
    InMux I__2865 (
            .O(N__24402),
            .I(N__24399));
    LocalMux I__2864 (
            .O(N__24399),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__2863 (
            .O(N__24396),
            .I(N__24393));
    LocalMux I__2862 (
            .O(N__24393),
            .I(N__24390));
    Span4Mux_v I__2861 (
            .O(N__24390),
            .I(N__24387));
    Odrv4 I__2860 (
            .O(N__24387),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__2859 (
            .O(N__24384),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__2858 (
            .O(N__24381),
            .I(N__24378));
    LocalMux I__2857 (
            .O(N__24378),
            .I(N__24375));
    Odrv12 I__2856 (
            .O(N__24375),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__2855 (
            .O(N__24372),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    CascadeMux I__2854 (
            .O(N__24369),
            .I(N__24366));
    InMux I__2853 (
            .O(N__24366),
            .I(N__24363));
    LocalMux I__2852 (
            .O(N__24363),
            .I(N__24360));
    Odrv4 I__2851 (
            .O(N__24360),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__2850 (
            .O(N__24357),
            .I(N__24354));
    LocalMux I__2849 (
            .O(N__24354),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__2848 (
            .O(N__24351),
            .I(bfn_8_14_0_));
    InMux I__2847 (
            .O(N__24348),
            .I(N__24345));
    LocalMux I__2846 (
            .O(N__24345),
            .I(N__24342));
    Odrv12 I__2845 (
            .O(N__24342),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__2844 (
            .O(N__24339),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__2843 (
            .O(N__24336),
            .I(N__24333));
    LocalMux I__2842 (
            .O(N__24333),
            .I(N__24330));
    Odrv12 I__2841 (
            .O(N__24330),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__2840 (
            .O(N__24327),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__2839 (
            .O(N__24324),
            .I(N__24321));
    LocalMux I__2838 (
            .O(N__24321),
            .I(N__24318));
    Span4Mux_h I__2837 (
            .O(N__24318),
            .I(N__24315));
    Odrv4 I__2836 (
            .O(N__24315),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__2835 (
            .O(N__24312),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__2834 (
            .O(N__24309),
            .I(N__24306));
    LocalMux I__2833 (
            .O(N__24306),
            .I(N__24303));
    Odrv12 I__2832 (
            .O(N__24303),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__2831 (
            .O(N__24300),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__2830 (
            .O(N__24297),
            .I(N__24294));
    LocalMux I__2829 (
            .O(N__24294),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__2828 (
            .O(N__24291),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__2827 (
            .O(N__24288),
            .I(N__24285));
    LocalMux I__2826 (
            .O(N__24285),
            .I(N__24282));
    Span4Mux_h I__2825 (
            .O(N__24282),
            .I(N__24279));
    Odrv4 I__2824 (
            .O(N__24279),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__2823 (
            .O(N__24276),
            .I(N__24273));
    LocalMux I__2822 (
            .O(N__24273),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__2821 (
            .O(N__24270),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__2820 (
            .O(N__24267),
            .I(N__24264));
    LocalMux I__2819 (
            .O(N__24264),
            .I(N__24261));
    Span4Mux_h I__2818 (
            .O(N__24261),
            .I(N__24258));
    Odrv4 I__2817 (
            .O(N__24258),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__2816 (
            .O(N__24255),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__2815 (
            .O(N__24252),
            .I(N__24249));
    LocalMux I__2814 (
            .O(N__24249),
            .I(N__24246));
    Odrv12 I__2813 (
            .O(N__24246),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__2812 (
            .O(N__24243),
            .I(bfn_8_13_0_));
    InMux I__2811 (
            .O(N__24240),
            .I(N__24237));
    LocalMux I__2810 (
            .O(N__24237),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__2809 (
            .O(N__24234),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__2808 (
            .O(N__24231),
            .I(N__24228));
    LocalMux I__2807 (
            .O(N__24228),
            .I(N__24225));
    Odrv4 I__2806 (
            .O(N__24225),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__2805 (
            .O(N__24222),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__2804 (
            .O(N__24219),
            .I(N__24216));
    LocalMux I__2803 (
            .O(N__24216),
            .I(N__24213));
    Span4Mux_v I__2802 (
            .O(N__24213),
            .I(N__24210));
    Odrv4 I__2801 (
            .O(N__24210),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__2800 (
            .O(N__24207),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__2799 (
            .O(N__24204),
            .I(N__24201));
    LocalMux I__2798 (
            .O(N__24201),
            .I(N__24198));
    Odrv4 I__2797 (
            .O(N__24198),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__2796 (
            .O(N__24195),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__2795 (
            .O(N__24192),
            .I(N__24189));
    LocalMux I__2794 (
            .O(N__24189),
            .I(N__24186));
    Odrv12 I__2793 (
            .O(N__24186),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__2792 (
            .O(N__24183),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__2791 (
            .O(N__24180),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    InMux I__2790 (
            .O(N__24177),
            .I(N__24174));
    LocalMux I__2789 (
            .O(N__24174),
            .I(N__24171));
    Span4Mux_v I__2788 (
            .O(N__24171),
            .I(N__24168));
    Odrv4 I__2787 (
            .O(N__24168),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__2786 (
            .O(N__24165),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__2785 (
            .O(N__24162),
            .I(N__24159));
    LocalMux I__2784 (
            .O(N__24159),
            .I(N__24156));
    Span4Mux_v I__2783 (
            .O(N__24156),
            .I(N__24153));
    Odrv4 I__2782 (
            .O(N__24153),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__2781 (
            .O(N__24150),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__2780 (
            .O(N__24147),
            .I(N__24144));
    LocalMux I__2779 (
            .O(N__24144),
            .I(N__24141));
    Odrv12 I__2778 (
            .O(N__24141),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__2777 (
            .O(N__24138),
            .I(bfn_8_12_0_));
    InMux I__2776 (
            .O(N__24135),
            .I(N__24132));
    LocalMux I__2775 (
            .O(N__24132),
            .I(N__24129));
    Odrv12 I__2774 (
            .O(N__24129),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__2773 (
            .O(N__24126),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__2772 (
            .O(N__24123),
            .I(N__24120));
    LocalMux I__2771 (
            .O(N__24120),
            .I(N__24117));
    Odrv12 I__2770 (
            .O(N__24117),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__2769 (
            .O(N__24114),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__2768 (
            .O(N__24111),
            .I(N__24108));
    LocalMux I__2767 (
            .O(N__24108),
            .I(N__24105));
    Odrv12 I__2766 (
            .O(N__24105),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__2765 (
            .O(N__24102),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__2764 (
            .O(N__24099),
            .I(N__24096));
    LocalMux I__2763 (
            .O(N__24096),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__2762 (
            .O(N__24093),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    CascadeMux I__2761 (
            .O(N__24090),
            .I(N__24087));
    InMux I__2760 (
            .O(N__24087),
            .I(N__24084));
    LocalMux I__2759 (
            .O(N__24084),
            .I(N__24081));
    Span4Mux_v I__2758 (
            .O(N__24081),
            .I(N__24078));
    Odrv4 I__2757 (
            .O(N__24078),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__2756 (
            .O(N__24075),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__2755 (
            .O(N__24072),
            .I(N__24063));
    InMux I__2754 (
            .O(N__24071),
            .I(N__24063));
    InMux I__2753 (
            .O(N__24070),
            .I(N__24063));
    LocalMux I__2752 (
            .O(N__24063),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    CascadeMux I__2751 (
            .O(N__24060),
            .I(N__24055));
    CascadeMux I__2750 (
            .O(N__24059),
            .I(N__24052));
    CascadeMux I__2749 (
            .O(N__24058),
            .I(N__24049));
    InMux I__2748 (
            .O(N__24055),
            .I(N__24042));
    InMux I__2747 (
            .O(N__24052),
            .I(N__24042));
    InMux I__2746 (
            .O(N__24049),
            .I(N__24042));
    LocalMux I__2745 (
            .O(N__24042),
            .I(\phase_controller_inst2.start_flagZ0 ));
    InMux I__2744 (
            .O(N__24039),
            .I(N__24036));
    LocalMux I__2743 (
            .O(N__24036),
            .I(\phase_controller_inst2.state_ns_0_0_1 ));
    InMux I__2742 (
            .O(N__24033),
            .I(N__24030));
    LocalMux I__2741 (
            .O(N__24030),
            .I(N__24027));
    Span4Mux_v I__2740 (
            .O(N__24027),
            .I(N__24024));
    Odrv4 I__2739 (
            .O(N__24024),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__2738 (
            .O(N__24021),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    InMux I__2737 (
            .O(N__24018),
            .I(N__24015));
    LocalMux I__2736 (
            .O(N__24015),
            .I(N__24012));
    Span4Mux_v I__2735 (
            .O(N__24012),
            .I(N__24009));
    Odrv4 I__2734 (
            .O(N__24009),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__2733 (
            .O(N__24006),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__2732 (
            .O(N__24003),
            .I(N__24000));
    LocalMux I__2731 (
            .O(N__24000),
            .I(N__23997));
    Span4Mux_v I__2730 (
            .O(N__23997),
            .I(N__23994));
    Odrv4 I__2729 (
            .O(N__23994),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__2728 (
            .O(N__23991),
            .I(N__23987));
    InMux I__2727 (
            .O(N__23990),
            .I(N__23984));
    LocalMux I__2726 (
            .O(N__23987),
            .I(N__23981));
    LocalMux I__2725 (
            .O(N__23984),
            .I(N__23978));
    Span4Mux_v I__2724 (
            .O(N__23981),
            .I(N__23975));
    Span4Mux_v I__2723 (
            .O(N__23978),
            .I(N__23972));
    Span4Mux_v I__2722 (
            .O(N__23975),
            .I(N__23969));
    Span4Mux_h I__2721 (
            .O(N__23972),
            .I(N__23966));
    Odrv4 I__2720 (
            .O(N__23969),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv4 I__2719 (
            .O(N__23966),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__2718 (
            .O(N__23961),
            .I(N__23958));
    LocalMux I__2717 (
            .O(N__23958),
            .I(N__23954));
    CascadeMux I__2716 (
            .O(N__23957),
            .I(N__23951));
    Span4Mux_v I__2715 (
            .O(N__23954),
            .I(N__23947));
    InMux I__2714 (
            .O(N__23951),
            .I(N__23942));
    InMux I__2713 (
            .O(N__23950),
            .I(N__23942));
    Sp12to4 I__2712 (
            .O(N__23947),
            .I(N__23937));
    LocalMux I__2711 (
            .O(N__23942),
            .I(N__23937));
    Span12Mux_h I__2710 (
            .O(N__23937),
            .I(N__23934));
    Odrv12 I__2709 (
            .O(N__23934),
            .I(il_max_comp2_c));
    InMux I__2708 (
            .O(N__23931),
            .I(N__23928));
    LocalMux I__2707 (
            .O(N__23928),
            .I(N__23925));
    Span4Mux_h I__2706 (
            .O(N__23925),
            .I(N__23922));
    Span4Mux_v I__2705 (
            .O(N__23922),
            .I(N__23919));
    Odrv4 I__2704 (
            .O(N__23919),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__2703 (
            .O(N__23916),
            .I(N__23912));
    InMux I__2702 (
            .O(N__23915),
            .I(N__23909));
    LocalMux I__2701 (
            .O(N__23912),
            .I(N__23906));
    LocalMux I__2700 (
            .O(N__23909),
            .I(N__23903));
    Span4Mux_v I__2699 (
            .O(N__23906),
            .I(N__23900));
    Span4Mux_s1_h I__2698 (
            .O(N__23903),
            .I(N__23897));
    Span4Mux_v I__2697 (
            .O(N__23900),
            .I(N__23894));
    Span4Mux_h I__2696 (
            .O(N__23897),
            .I(N__23891));
    Odrv4 I__2695 (
            .O(N__23894),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__2694 (
            .O(N__23891),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__2693 (
            .O(N__23886),
            .I(N__23883));
    LocalMux I__2692 (
            .O(N__23883),
            .I(N__23879));
    InMux I__2691 (
            .O(N__23882),
            .I(N__23876));
    Span4Mux_v I__2690 (
            .O(N__23879),
            .I(N__23873));
    LocalMux I__2689 (
            .O(N__23876),
            .I(N__23870));
    Span4Mux_v I__2688 (
            .O(N__23873),
            .I(N__23865));
    Span4Mux_s3_h I__2687 (
            .O(N__23870),
            .I(N__23865));
    Odrv4 I__2686 (
            .O(N__23865),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__2685 (
            .O(N__23862),
            .I(N__23859));
    LocalMux I__2684 (
            .O(N__23859),
            .I(N__23856));
    Span4Mux_v I__2683 (
            .O(N__23856),
            .I(N__23852));
    InMux I__2682 (
            .O(N__23855),
            .I(N__23849));
    Span4Mux_v I__2681 (
            .O(N__23852),
            .I(N__23846));
    LocalMux I__2680 (
            .O(N__23849),
            .I(N__23843));
    Odrv4 I__2679 (
            .O(N__23846),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv12 I__2678 (
            .O(N__23843),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__2677 (
            .O(N__23838),
            .I(N__23834));
    InMux I__2676 (
            .O(N__23837),
            .I(N__23831));
    LocalMux I__2675 (
            .O(N__23834),
            .I(N__23828));
    LocalMux I__2674 (
            .O(N__23831),
            .I(N__23825));
    Span4Mux_h I__2673 (
            .O(N__23828),
            .I(N__23822));
    Span4Mux_v I__2672 (
            .O(N__23825),
            .I(N__23819));
    Span4Mux_v I__2671 (
            .O(N__23822),
            .I(N__23816));
    Span4Mux_h I__2670 (
            .O(N__23819),
            .I(N__23813));
    Odrv4 I__2669 (
            .O(N__23816),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv4 I__2668 (
            .O(N__23813),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__2667 (
            .O(N__23808),
            .I(N__23804));
    InMux I__2666 (
            .O(N__23807),
            .I(N__23801));
    LocalMux I__2665 (
            .O(N__23804),
            .I(N__23798));
    LocalMux I__2664 (
            .O(N__23801),
            .I(N__23795));
    Span4Mux_h I__2663 (
            .O(N__23798),
            .I(N__23792));
    Span4Mux_v I__2662 (
            .O(N__23795),
            .I(N__23789));
    Span4Mux_v I__2661 (
            .O(N__23792),
            .I(N__23786));
    Span4Mux_h I__2660 (
            .O(N__23789),
            .I(N__23783));
    Odrv4 I__2659 (
            .O(N__23786),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    Odrv4 I__2658 (
            .O(N__23783),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__2657 (
            .O(N__23778),
            .I(N__23774));
    InMux I__2656 (
            .O(N__23777),
            .I(N__23771));
    LocalMux I__2655 (
            .O(N__23774),
            .I(N__23768));
    LocalMux I__2654 (
            .O(N__23771),
            .I(N__23765));
    Span4Mux_v I__2653 (
            .O(N__23768),
            .I(N__23762));
    Span4Mux_v I__2652 (
            .O(N__23765),
            .I(N__23759));
    Span4Mux_v I__2651 (
            .O(N__23762),
            .I(N__23756));
    Span4Mux_h I__2650 (
            .O(N__23759),
            .I(N__23753));
    Odrv4 I__2649 (
            .O(N__23756),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv4 I__2648 (
            .O(N__23753),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__2647 (
            .O(N__23748),
            .I(N__23745));
    LocalMux I__2646 (
            .O(N__23745),
            .I(N__23742));
    Span4Mux_v I__2645 (
            .O(N__23742),
            .I(N__23738));
    InMux I__2644 (
            .O(N__23741),
            .I(N__23735));
    Sp12to4 I__2643 (
            .O(N__23738),
            .I(N__23730));
    LocalMux I__2642 (
            .O(N__23735),
            .I(N__23730));
    Span12Mux_s5_h I__2641 (
            .O(N__23730),
            .I(N__23727));
    Odrv12 I__2640 (
            .O(N__23727),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__2639 (
            .O(N__23724),
            .I(N__23720));
    InMux I__2638 (
            .O(N__23723),
            .I(N__23717));
    LocalMux I__2637 (
            .O(N__23720),
            .I(N__23714));
    LocalMux I__2636 (
            .O(N__23717),
            .I(N__23711));
    Span4Mux_h I__2635 (
            .O(N__23714),
            .I(N__23708));
    Span12Mux_s5_h I__2634 (
            .O(N__23711),
            .I(N__23705));
    Odrv4 I__2633 (
            .O(N__23708),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    Odrv12 I__2632 (
            .O(N__23705),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__2631 (
            .O(N__23700),
            .I(N__23697));
    LocalMux I__2630 (
            .O(N__23697),
            .I(N__23694));
    Span4Mux_h I__2629 (
            .O(N__23694),
            .I(N__23691));
    Odrv4 I__2628 (
            .O(N__23691),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__2627 (
            .O(N__23688),
            .I(N__23685));
    LocalMux I__2626 (
            .O(N__23685),
            .I(N__23682));
    Span4Mux_v I__2625 (
            .O(N__23682),
            .I(N__23679));
    Span4Mux_h I__2624 (
            .O(N__23679),
            .I(N__23676));
    Odrv4 I__2623 (
            .O(N__23676),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__2622 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__2621 (
            .O(N__23670),
            .I(N__23666));
    InMux I__2620 (
            .O(N__23669),
            .I(N__23663));
    Span4Mux_v I__2619 (
            .O(N__23666),
            .I(N__23658));
    LocalMux I__2618 (
            .O(N__23663),
            .I(N__23658));
    Span4Mux_h I__2617 (
            .O(N__23658),
            .I(N__23655));
    Span4Mux_v I__2616 (
            .O(N__23655),
            .I(N__23652));
    Odrv4 I__2615 (
            .O(N__23652),
            .I(\current_shift_inst.control_input_axb_0 ));
    InMux I__2614 (
            .O(N__23649),
            .I(N__23646));
    LocalMux I__2613 (
            .O(N__23646),
            .I(N__23643));
    Span4Mux_h I__2612 (
            .O(N__23643),
            .I(N__23640));
    Span4Mux_v I__2611 (
            .O(N__23640),
            .I(N__23637));
    Odrv4 I__2610 (
            .O(N__23637),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__2609 (
            .O(N__23634),
            .I(N__23631));
    LocalMux I__2608 (
            .O(N__23631),
            .I(N__23628));
    Span12Mux_s7_h I__2607 (
            .O(N__23628),
            .I(N__23625));
    Odrv12 I__2606 (
            .O(N__23625),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__2605 (
            .O(N__23622),
            .I(N__23619));
    LocalMux I__2604 (
            .O(N__23619),
            .I(N__23615));
    InMux I__2603 (
            .O(N__23618),
            .I(N__23612));
    Span4Mux_s1_h I__2602 (
            .O(N__23615),
            .I(N__23609));
    LocalMux I__2601 (
            .O(N__23612),
            .I(N__23606));
    Span4Mux_h I__2600 (
            .O(N__23609),
            .I(N__23603));
    Odrv4 I__2599 (
            .O(N__23606),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__2598 (
            .O(N__23603),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__2597 (
            .O(N__23598),
            .I(N__23595));
    LocalMux I__2596 (
            .O(N__23595),
            .I(N__23592));
    Span4Mux_h I__2595 (
            .O(N__23592),
            .I(N__23589));
    Odrv4 I__2594 (
            .O(N__23589),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__2593 (
            .O(N__23586),
            .I(N__23583));
    LocalMux I__2592 (
            .O(N__23583),
            .I(N__23580));
    Span4Mux_h I__2591 (
            .O(N__23580),
            .I(N__23577));
    Odrv4 I__2590 (
            .O(N__23577),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__2589 (
            .O(N__23574),
            .I(N__23571));
    LocalMux I__2588 (
            .O(N__23571),
            .I(N__23568));
    Span4Mux_h I__2587 (
            .O(N__23568),
            .I(N__23565));
    Odrv4 I__2586 (
            .O(N__23565),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__2585 (
            .O(N__23562),
            .I(N__23559));
    LocalMux I__2584 (
            .O(N__23559),
            .I(N__23556));
    Odrv12 I__2583 (
            .O(N__23556),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__2582 (
            .O(N__23553),
            .I(N__23550));
    LocalMux I__2581 (
            .O(N__23550),
            .I(N__23547));
    Span4Mux_h I__2580 (
            .O(N__23547),
            .I(N__23544));
    Odrv4 I__2579 (
            .O(N__23544),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__2578 (
            .O(N__23541),
            .I(N__23538));
    LocalMux I__2577 (
            .O(N__23538),
            .I(N__23535));
    Span4Mux_h I__2576 (
            .O(N__23535),
            .I(N__23532));
    Odrv4 I__2575 (
            .O(N__23532),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__2574 (
            .O(N__23529),
            .I(N__23526));
    LocalMux I__2573 (
            .O(N__23526),
            .I(N__23523));
    Span4Mux_h I__2572 (
            .O(N__23523),
            .I(N__23520));
    Odrv4 I__2571 (
            .O(N__23520),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__2570 (
            .O(N__23517),
            .I(N__23513));
    InMux I__2569 (
            .O(N__23516),
            .I(N__23510));
    LocalMux I__2568 (
            .O(N__23513),
            .I(N__23507));
    LocalMux I__2567 (
            .O(N__23510),
            .I(N__23504));
    Span4Mux_s1_h I__2566 (
            .O(N__23507),
            .I(N__23501));
    Span4Mux_v I__2565 (
            .O(N__23504),
            .I(N__23498));
    Span4Mux_h I__2564 (
            .O(N__23501),
            .I(N__23495));
    Odrv4 I__2563 (
            .O(N__23498),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__2562 (
            .O(N__23495),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__2561 (
            .O(N__23490),
            .I(N__23486));
    InMux I__2560 (
            .O(N__23489),
            .I(N__23483));
    LocalMux I__2559 (
            .O(N__23486),
            .I(N__23480));
    LocalMux I__2558 (
            .O(N__23483),
            .I(N__23477));
    Span4Mux_v I__2557 (
            .O(N__23480),
            .I(N__23474));
    Span4Mux_v I__2556 (
            .O(N__23477),
            .I(N__23471));
    Span4Mux_h I__2555 (
            .O(N__23474),
            .I(N__23468));
    Odrv4 I__2554 (
            .O(N__23471),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    Odrv4 I__2553 (
            .O(N__23468),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__2552 (
            .O(N__23463),
            .I(N__23460));
    LocalMux I__2551 (
            .O(N__23460),
            .I(N__23456));
    InMux I__2550 (
            .O(N__23459),
            .I(N__23453));
    Span4Mux_v I__2549 (
            .O(N__23456),
            .I(N__23450));
    LocalMux I__2548 (
            .O(N__23453),
            .I(N__23447));
    Span4Mux_h I__2547 (
            .O(N__23450),
            .I(N__23444));
    Odrv12 I__2546 (
            .O(N__23447),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv4 I__2545 (
            .O(N__23444),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__2544 (
            .O(N__23439),
            .I(N__23436));
    LocalMux I__2543 (
            .O(N__23436),
            .I(N__23432));
    InMux I__2542 (
            .O(N__23435),
            .I(N__23429));
    Span4Mux_v I__2541 (
            .O(N__23432),
            .I(N__23426));
    LocalMux I__2540 (
            .O(N__23429),
            .I(N__23423));
    Span4Mux_h I__2539 (
            .O(N__23426),
            .I(N__23420));
    Odrv12 I__2538 (
            .O(N__23423),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv4 I__2537 (
            .O(N__23420),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__2536 (
            .O(N__23415),
            .I(N__23412));
    LocalMux I__2535 (
            .O(N__23412),
            .I(N__23409));
    Odrv12 I__2534 (
            .O(N__23409),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__2533 (
            .O(N__23406),
            .I(N__23403));
    LocalMux I__2532 (
            .O(N__23403),
            .I(N__23400));
    Span4Mux_s1_h I__2531 (
            .O(N__23400),
            .I(N__23396));
    InMux I__2530 (
            .O(N__23399),
            .I(N__23393));
    Span4Mux_v I__2529 (
            .O(N__23396),
            .I(N__23390));
    LocalMux I__2528 (
            .O(N__23393),
            .I(N__23387));
    Span4Mux_h I__2527 (
            .O(N__23390),
            .I(N__23384));
    Odrv12 I__2526 (
            .O(N__23387),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv4 I__2525 (
            .O(N__23384),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__2524 (
            .O(N__23379),
            .I(N__23375));
    InMux I__2523 (
            .O(N__23378),
            .I(N__23372));
    LocalMux I__2522 (
            .O(N__23375),
            .I(N__23369));
    LocalMux I__2521 (
            .O(N__23372),
            .I(N__23366));
    Span12Mux_v I__2520 (
            .O(N__23369),
            .I(N__23363));
    Odrv12 I__2519 (
            .O(N__23366),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv12 I__2518 (
            .O(N__23363),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__2517 (
            .O(N__23358),
            .I(N__23355));
    LocalMux I__2516 (
            .O(N__23355),
            .I(N__23351));
    InMux I__2515 (
            .O(N__23354),
            .I(N__23348));
    Span4Mux_v I__2514 (
            .O(N__23351),
            .I(N__23345));
    LocalMux I__2513 (
            .O(N__23348),
            .I(N__23342));
    Span4Mux_v I__2512 (
            .O(N__23345),
            .I(N__23339));
    Span12Mux_s10_v I__2511 (
            .O(N__23342),
            .I(N__23336));
    Span4Mux_h I__2510 (
            .O(N__23339),
            .I(N__23333));
    Odrv12 I__2509 (
            .O(N__23336),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    Odrv4 I__2508 (
            .O(N__23333),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    ClkMux I__2507 (
            .O(N__23328),
            .I(N__23325));
    GlobalMux I__2506 (
            .O(N__23325),
            .I(N__23322));
    gio2CtrlBuf I__2505 (
            .O(N__23322),
            .I(delay_hc_input_c_g));
    InMux I__2504 (
            .O(N__23319),
            .I(N__23315));
    InMux I__2503 (
            .O(N__23318),
            .I(N__23312));
    LocalMux I__2502 (
            .O(N__23315),
            .I(N__23309));
    LocalMux I__2501 (
            .O(N__23312),
            .I(N__23306));
    Span4Mux_s2_h I__2500 (
            .O(N__23309),
            .I(N__23303));
    Odrv4 I__2499 (
            .O(N__23306),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__2498 (
            .O(N__23303),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__2497 (
            .O(N__23298),
            .I(N__23294));
    InMux I__2496 (
            .O(N__23297),
            .I(N__23291));
    LocalMux I__2495 (
            .O(N__23294),
            .I(N__23288));
    LocalMux I__2494 (
            .O(N__23291),
            .I(N__23285));
    Odrv12 I__2493 (
            .O(N__23288),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__2492 (
            .O(N__23285),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__2491 (
            .O(N__23280),
            .I(N__23276));
    InMux I__2490 (
            .O(N__23279),
            .I(N__23273));
    LocalMux I__2489 (
            .O(N__23276),
            .I(N__23270));
    LocalMux I__2488 (
            .O(N__23273),
            .I(N__23267));
    Span4Mux_s3_h I__2487 (
            .O(N__23270),
            .I(N__23264));
    Odrv12 I__2486 (
            .O(N__23267),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__2485 (
            .O(N__23264),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__2484 (
            .O(N__23259),
            .I(N__23256));
    LocalMux I__2483 (
            .O(N__23256),
            .I(N__23252));
    InMux I__2482 (
            .O(N__23255),
            .I(N__23249));
    Span4Mux_v I__2481 (
            .O(N__23252),
            .I(N__23246));
    LocalMux I__2480 (
            .O(N__23249),
            .I(N__23243));
    Span4Mux_h I__2479 (
            .O(N__23246),
            .I(N__23240));
    Odrv4 I__2478 (
            .O(N__23243),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    Odrv4 I__2477 (
            .O(N__23240),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__2476 (
            .O(N__23235),
            .I(N__23232));
    LocalMux I__2475 (
            .O(N__23232),
            .I(N__23228));
    InMux I__2474 (
            .O(N__23231),
            .I(N__23225));
    Span4Mux_v I__2473 (
            .O(N__23228),
            .I(N__23222));
    LocalMux I__2472 (
            .O(N__23225),
            .I(N__23219));
    Span4Mux_h I__2471 (
            .O(N__23222),
            .I(N__23216));
    Odrv4 I__2470 (
            .O(N__23219),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    Odrv4 I__2469 (
            .O(N__23216),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__2468 (
            .O(N__23211),
            .I(N__23208));
    LocalMux I__2467 (
            .O(N__23208),
            .I(N__23204));
    InMux I__2466 (
            .O(N__23207),
            .I(N__23201));
    Span4Mux_v I__2465 (
            .O(N__23204),
            .I(N__23198));
    LocalMux I__2464 (
            .O(N__23201),
            .I(N__23195));
    Span4Mux_h I__2463 (
            .O(N__23198),
            .I(N__23192));
    Odrv4 I__2462 (
            .O(N__23195),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    Odrv4 I__2461 (
            .O(N__23192),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__2460 (
            .O(N__23187),
            .I(N__23184));
    LocalMux I__2459 (
            .O(N__23184),
            .I(N__23180));
    InMux I__2458 (
            .O(N__23183),
            .I(N__23177));
    Span4Mux_v I__2457 (
            .O(N__23180),
            .I(N__23174));
    LocalMux I__2456 (
            .O(N__23177),
            .I(N__23171));
    Span4Mux_h I__2455 (
            .O(N__23174),
            .I(N__23168));
    Odrv12 I__2454 (
            .O(N__23171),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv4 I__2453 (
            .O(N__23168),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__2452 (
            .O(N__23163),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__2451 (
            .O(N__23160),
            .I(N__23157));
    LocalMux I__2450 (
            .O(N__23157),
            .I(N__23154));
    Odrv4 I__2449 (
            .O(N__23154),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__2448 (
            .O(N__23151),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__2447 (
            .O(N__23148),
            .I(N__23145));
    LocalMux I__2446 (
            .O(N__23145),
            .I(N__23142));
    Odrv4 I__2445 (
            .O(N__23142),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__2444 (
            .O(N__23139),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__2443 (
            .O(N__23136),
            .I(N__23133));
    LocalMux I__2442 (
            .O(N__23133),
            .I(N__23130));
    Odrv12 I__2441 (
            .O(N__23130),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__2440 (
            .O(N__23127),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__2439 (
            .O(N__23124),
            .I(N__23121));
    LocalMux I__2438 (
            .O(N__23121),
            .I(N__23118));
    Odrv12 I__2437 (
            .O(N__23118),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__2436 (
            .O(N__23115),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__2435 (
            .O(N__23112),
            .I(N__23109));
    LocalMux I__2434 (
            .O(N__23109),
            .I(N__23106));
    Odrv4 I__2433 (
            .O(N__23106),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    InMux I__2432 (
            .O(N__23103),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__2431 (
            .O(N__23100),
            .I(N__23097));
    LocalMux I__2430 (
            .O(N__23097),
            .I(N__23094));
    Odrv4 I__2429 (
            .O(N__23094),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__2428 (
            .O(N__23091),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__2427 (
            .O(N__23088),
            .I(N__23084));
    InMux I__2426 (
            .O(N__23087),
            .I(N__23081));
    LocalMux I__2425 (
            .O(N__23084),
            .I(N__23078));
    LocalMux I__2424 (
            .O(N__23081),
            .I(N__23075));
    Span4Mux_s1_h I__2423 (
            .O(N__23078),
            .I(N__23072));
    Span4Mux_v I__2422 (
            .O(N__23075),
            .I(N__23067));
    Span4Mux_h I__2421 (
            .O(N__23072),
            .I(N__23067));
    Odrv4 I__2420 (
            .O(N__23067),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__2419 (
            .O(N__23064),
            .I(N__23061));
    LocalMux I__2418 (
            .O(N__23061),
            .I(N__23057));
    InMux I__2417 (
            .O(N__23060),
            .I(N__23054));
    Span4Mux_v I__2416 (
            .O(N__23057),
            .I(N__23051));
    LocalMux I__2415 (
            .O(N__23054),
            .I(N__23048));
    Span4Mux_h I__2414 (
            .O(N__23051),
            .I(N__23045));
    Odrv4 I__2413 (
            .O(N__23048),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__2412 (
            .O(N__23045),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__2411 (
            .O(N__23040),
            .I(N__23037));
    LocalMux I__2410 (
            .O(N__23037),
            .I(N__23034));
    Odrv4 I__2409 (
            .O(N__23034),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__2408 (
            .O(N__23031),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__2407 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__2406 (
            .O(N__23025),
            .I(N__23022));
    Odrv4 I__2405 (
            .O(N__23022),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__2404 (
            .O(N__23019),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__2403 (
            .O(N__23016),
            .I(N__23013));
    LocalMux I__2402 (
            .O(N__23013),
            .I(N__23010));
    Odrv4 I__2401 (
            .O(N__23010),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__2400 (
            .O(N__23007),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__2399 (
            .O(N__23004),
            .I(N__23001));
    LocalMux I__2398 (
            .O(N__23001),
            .I(N__22998));
    Odrv12 I__2397 (
            .O(N__22998),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__2396 (
            .O(N__22995),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__2395 (
            .O(N__22992),
            .I(N__22989));
    LocalMux I__2394 (
            .O(N__22989),
            .I(N__22986));
    Odrv12 I__2393 (
            .O(N__22986),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__2392 (
            .O(N__22983),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__2391 (
            .O(N__22980),
            .I(N__22977));
    LocalMux I__2390 (
            .O(N__22977),
            .I(N__22974));
    Odrv12 I__2389 (
            .O(N__22974),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__2388 (
            .O(N__22971),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    CascadeMux I__2387 (
            .O(N__22968),
            .I(N__22965));
    InMux I__2386 (
            .O(N__22965),
            .I(N__22962));
    LocalMux I__2385 (
            .O(N__22962),
            .I(N__22959));
    Odrv4 I__2384 (
            .O(N__22959),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__2383 (
            .O(N__22956),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__2382 (
            .O(N__22953),
            .I(N__22950));
    LocalMux I__2381 (
            .O(N__22950),
            .I(N__22947));
    Odrv4 I__2380 (
            .O(N__22947),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__2379 (
            .O(N__22944),
            .I(bfn_5_14_0_));
    InMux I__2378 (
            .O(N__22941),
            .I(N__22938));
    LocalMux I__2377 (
            .O(N__22938),
            .I(N__22935));
    Odrv4 I__2376 (
            .O(N__22935),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__2375 (
            .O(N__22932),
            .I(N__22929));
    LocalMux I__2374 (
            .O(N__22929),
            .I(N__22926));
    Odrv4 I__2373 (
            .O(N__22926),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__2372 (
            .O(N__22923),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__2371 (
            .O(N__22920),
            .I(N__22917));
    LocalMux I__2370 (
            .O(N__22917),
            .I(N__22914));
    Odrv4 I__2369 (
            .O(N__22914),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__2368 (
            .O(N__22911),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    CascadeMux I__2367 (
            .O(N__22908),
            .I(N__22905));
    InMux I__2366 (
            .O(N__22905),
            .I(N__22902));
    LocalMux I__2365 (
            .O(N__22902),
            .I(N__22899));
    Odrv4 I__2364 (
            .O(N__22899),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__2363 (
            .O(N__22896),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__2362 (
            .O(N__22893),
            .I(N__22890));
    LocalMux I__2361 (
            .O(N__22890),
            .I(N__22887));
    Odrv12 I__2360 (
            .O(N__22887),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__2359 (
            .O(N__22884),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__2358 (
            .O(N__22881),
            .I(N__22878));
    LocalMux I__2357 (
            .O(N__22878),
            .I(N__22875));
    Odrv12 I__2356 (
            .O(N__22875),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__2355 (
            .O(N__22872),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__2354 (
            .O(N__22869),
            .I(N__22866));
    LocalMux I__2353 (
            .O(N__22866),
            .I(N__22863));
    Odrv12 I__2352 (
            .O(N__22863),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__2351 (
            .O(N__22860),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__2350 (
            .O(N__22857),
            .I(N__22854));
    LocalMux I__2349 (
            .O(N__22854),
            .I(N__22851));
    Odrv4 I__2348 (
            .O(N__22851),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__2347 (
            .O(N__22848),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__2346 (
            .O(N__22845),
            .I(N__22842));
    LocalMux I__2345 (
            .O(N__22842),
            .I(N__22839));
    Odrv4 I__2344 (
            .O(N__22839),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__2343 (
            .O(N__22836),
            .I(bfn_5_13_0_));
    InMux I__2342 (
            .O(N__22833),
            .I(N__22830));
    LocalMux I__2341 (
            .O(N__22830),
            .I(N__22827));
    Odrv4 I__2340 (
            .O(N__22827),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__2339 (
            .O(N__22824),
            .I(N__22821));
    LocalMux I__2338 (
            .O(N__22821),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__2337 (
            .O(N__22818),
            .I(N__22815));
    LocalMux I__2336 (
            .O(N__22815),
            .I(N__22812));
    Odrv4 I__2335 (
            .O(N__22812),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__2334 (
            .O(N__22809),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    CascadeMux I__2333 (
            .O(N__22806),
            .I(N__22803));
    InMux I__2332 (
            .O(N__22803),
            .I(N__22800));
    LocalMux I__2331 (
            .O(N__22800),
            .I(N__22797));
    Odrv4 I__2330 (
            .O(N__22797),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__2329 (
            .O(N__22794),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__2328 (
            .O(N__22791),
            .I(N__22788));
    LocalMux I__2327 (
            .O(N__22788),
            .I(N__22785));
    Odrv4 I__2326 (
            .O(N__22785),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__2325 (
            .O(N__22782),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__2324 (
            .O(N__22779),
            .I(N__22776));
    LocalMux I__2323 (
            .O(N__22776),
            .I(N__22773));
    Odrv12 I__2322 (
            .O(N__22773),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__2321 (
            .O(N__22770),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__2320 (
            .O(N__22767),
            .I(N__22764));
    LocalMux I__2319 (
            .O(N__22764),
            .I(N__22761));
    Odrv12 I__2318 (
            .O(N__22761),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__2317 (
            .O(N__22758),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__2316 (
            .O(N__22755),
            .I(N__22752));
    LocalMux I__2315 (
            .O(N__22752),
            .I(N__22749));
    Odrv4 I__2314 (
            .O(N__22749),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__2313 (
            .O(N__22746),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__2312 (
            .O(N__22743),
            .I(N__22740));
    LocalMux I__2311 (
            .O(N__22740),
            .I(N__22737));
    Odrv12 I__2310 (
            .O(N__22737),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__2309 (
            .O(N__22734),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__2308 (
            .O(N__22731),
            .I(N__22728));
    LocalMux I__2307 (
            .O(N__22728),
            .I(N__22725));
    Odrv4 I__2306 (
            .O(N__22725),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__2305 (
            .O(N__22722),
            .I(bfn_5_12_0_));
    InMux I__2304 (
            .O(N__22719),
            .I(N__22716));
    LocalMux I__2303 (
            .O(N__22716),
            .I(\current_shift_inst.control_input_axb_23 ));
    InMux I__2302 (
            .O(N__22713),
            .I(N__22710));
    LocalMux I__2301 (
            .O(N__22710),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__2300 (
            .O(N__22707),
            .I(N__22704));
    LocalMux I__2299 (
            .O(N__22704),
            .I(N__22701));
    Span4Mux_h I__2298 (
            .O(N__22701),
            .I(N__22698));
    Odrv4 I__2297 (
            .O(N__22698),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__2296 (
            .O(N__22695),
            .I(N__22692));
    LocalMux I__2295 (
            .O(N__22692),
            .I(\current_shift_inst.control_input_axb_29 ));
    CascadeMux I__2294 (
            .O(N__22689),
            .I(\current_shift_inst.PI_CTRL.N_46_16_cascade_ ));
    InMux I__2293 (
            .O(N__22686),
            .I(N__22683));
    LocalMux I__2292 (
            .O(N__22683),
            .I(N__22680));
    Odrv12 I__2291 (
            .O(N__22680),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ));
    InMux I__2290 (
            .O(N__22677),
            .I(N__22674));
    LocalMux I__2289 (
            .O(N__22674),
            .I(N__22670));
    InMux I__2288 (
            .O(N__22673),
            .I(N__22667));
    Span4Mux_v I__2287 (
            .O(N__22670),
            .I(N__22664));
    LocalMux I__2286 (
            .O(N__22667),
            .I(N__22661));
    Span4Mux_v I__2285 (
            .O(N__22664),
            .I(N__22656));
    Span4Mux_h I__2284 (
            .O(N__22661),
            .I(N__22656));
    Odrv4 I__2283 (
            .O(N__22656),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    CascadeMux I__2282 (
            .O(N__22653),
            .I(N__22643));
    CascadeMux I__2281 (
            .O(N__22652),
            .I(N__22640));
    CascadeMux I__2280 (
            .O(N__22651),
            .I(N__22637));
    CascadeMux I__2279 (
            .O(N__22650),
            .I(N__22634));
    CEMux I__2278 (
            .O(N__22649),
            .I(N__22629));
    InMux I__2277 (
            .O(N__22648),
            .I(N__22617));
    InMux I__2276 (
            .O(N__22647),
            .I(N__22614));
    InMux I__2275 (
            .O(N__22646),
            .I(N__22611));
    InMux I__2274 (
            .O(N__22643),
            .I(N__22598));
    InMux I__2273 (
            .O(N__22640),
            .I(N__22598));
    InMux I__2272 (
            .O(N__22637),
            .I(N__22598));
    InMux I__2271 (
            .O(N__22634),
            .I(N__22598));
    InMux I__2270 (
            .O(N__22633),
            .I(N__22598));
    InMux I__2269 (
            .O(N__22632),
            .I(N__22598));
    LocalMux I__2268 (
            .O(N__22629),
            .I(N__22592));
    InMux I__2267 (
            .O(N__22628),
            .I(N__22587));
    InMux I__2266 (
            .O(N__22627),
            .I(N__22587));
    InMux I__2265 (
            .O(N__22626),
            .I(N__22580));
    InMux I__2264 (
            .O(N__22625),
            .I(N__22580));
    InMux I__2263 (
            .O(N__22624),
            .I(N__22580));
    InMux I__2262 (
            .O(N__22623),
            .I(N__22573));
    InMux I__2261 (
            .O(N__22622),
            .I(N__22573));
    InMux I__2260 (
            .O(N__22621),
            .I(N__22573));
    InMux I__2259 (
            .O(N__22620),
            .I(N__22570));
    LocalMux I__2258 (
            .O(N__22617),
            .I(N__22567));
    LocalMux I__2257 (
            .O(N__22614),
            .I(N__22564));
    LocalMux I__2256 (
            .O(N__22611),
            .I(N__22559));
    LocalMux I__2255 (
            .O(N__22598),
            .I(N__22559));
    InMux I__2254 (
            .O(N__22597),
            .I(N__22545));
    InMux I__2253 (
            .O(N__22596),
            .I(N__22545));
    InMux I__2252 (
            .O(N__22595),
            .I(N__22542));
    Span4Mux_h I__2251 (
            .O(N__22592),
            .I(N__22533));
    LocalMux I__2250 (
            .O(N__22587),
            .I(N__22533));
    LocalMux I__2249 (
            .O(N__22580),
            .I(N__22533));
    LocalMux I__2248 (
            .O(N__22573),
            .I(N__22533));
    LocalMux I__2247 (
            .O(N__22570),
            .I(N__22528));
    Span4Mux_h I__2246 (
            .O(N__22567),
            .I(N__22528));
    Span4Mux_h I__2245 (
            .O(N__22564),
            .I(N__22523));
    Span4Mux_h I__2244 (
            .O(N__22559),
            .I(N__22523));
    InMux I__2243 (
            .O(N__22558),
            .I(N__22520));
    InMux I__2242 (
            .O(N__22557),
            .I(N__22511));
    InMux I__2241 (
            .O(N__22556),
            .I(N__22511));
    InMux I__2240 (
            .O(N__22555),
            .I(N__22511));
    InMux I__2239 (
            .O(N__22554),
            .I(N__22511));
    InMux I__2238 (
            .O(N__22553),
            .I(N__22502));
    InMux I__2237 (
            .O(N__22552),
            .I(N__22502));
    InMux I__2236 (
            .O(N__22551),
            .I(N__22502));
    InMux I__2235 (
            .O(N__22550),
            .I(N__22502));
    LocalMux I__2234 (
            .O(N__22545),
            .I(N__22499));
    LocalMux I__2233 (
            .O(N__22542),
            .I(N__22494));
    Span4Mux_v I__2232 (
            .O(N__22533),
            .I(N__22494));
    Span4Mux_v I__2231 (
            .O(N__22528),
            .I(N__22491));
    Span4Mux_v I__2230 (
            .O(N__22523),
            .I(N__22488));
    LocalMux I__2229 (
            .O(N__22520),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__2228 (
            .O(N__22511),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__2227 (
            .O(N__22502),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv12 I__2226 (
            .O(N__22499),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__2225 (
            .O(N__22494),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__2224 (
            .O(N__22491),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__2223 (
            .O(N__22488),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    InMux I__2222 (
            .O(N__22473),
            .I(N__22470));
    LocalMux I__2221 (
            .O(N__22470),
            .I(N__22467));
    Span4Mux_v I__2220 (
            .O(N__22467),
            .I(N__22464));
    Odrv4 I__2219 (
            .O(N__22464),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__2218 (
            .O(N__22461),
            .I(N__22458));
    LocalMux I__2217 (
            .O(N__22458),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__2216 (
            .O(N__22455),
            .I(N__22452));
    LocalMux I__2215 (
            .O(N__22452),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__2214 (
            .O(N__22449),
            .I(N__22446));
    LocalMux I__2213 (
            .O(N__22446),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__2212 (
            .O(N__22443),
            .I(N__22440));
    LocalMux I__2211 (
            .O(N__22440),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__2210 (
            .O(N__22437),
            .I(N__22434));
    LocalMux I__2209 (
            .O(N__22434),
            .I(\current_shift_inst.control_input_axb_20 ));
    InMux I__2208 (
            .O(N__22431),
            .I(N__22428));
    LocalMux I__2207 (
            .O(N__22428),
            .I(N__22425));
    Odrv12 I__2206 (
            .O(N__22425),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    InMux I__2205 (
            .O(N__22422),
            .I(N__22419));
    LocalMux I__2204 (
            .O(N__22419),
            .I(N__22416));
    Odrv4 I__2203 (
            .O(N__22416),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__2202 (
            .O(N__22413),
            .I(N__22410));
    LocalMux I__2201 (
            .O(N__22410),
            .I(\current_shift_inst.control_input_axb_27 ));
    InMux I__2200 (
            .O(N__22407),
            .I(N__22404));
    LocalMux I__2199 (
            .O(N__22404),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__2198 (
            .O(N__22401),
            .I(N__22398));
    LocalMux I__2197 (
            .O(N__22398),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__2196 (
            .O(N__22395),
            .I(N__22392));
    LocalMux I__2195 (
            .O(N__22392),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__2194 (
            .O(N__22389),
            .I(N__22386));
    LocalMux I__2193 (
            .O(N__22386),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    InMux I__2192 (
            .O(N__22383),
            .I(N__22380));
    LocalMux I__2191 (
            .O(N__22380),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__2190 (
            .O(N__22377),
            .I(N__22374));
    LocalMux I__2189 (
            .O(N__22374),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__2188 (
            .O(N__22371),
            .I(N__22368));
    LocalMux I__2187 (
            .O(N__22368),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__2186 (
            .O(N__22365),
            .I(N__22362));
    LocalMux I__2185 (
            .O(N__22362),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__2184 (
            .O(N__22359),
            .I(N__22356));
    LocalMux I__2183 (
            .O(N__22356),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__2182 (
            .O(N__22353),
            .I(N__22350));
    LocalMux I__2181 (
            .O(N__22350),
            .I(\current_shift_inst.control_input_axb_12 ));
    CascadeMux I__2180 (
            .O(N__22347),
            .I(N__22344));
    InMux I__2179 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__2178 (
            .O(N__22341),
            .I(N__22338));
    Odrv4 I__2177 (
            .O(N__22338),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__2176 (
            .O(N__22335),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ));
    InMux I__2175 (
            .O(N__22332),
            .I(N__22329));
    LocalMux I__2174 (
            .O(N__22329),
            .I(\current_shift_inst.PI_CTRL.N_77 ));
    CascadeMux I__2173 (
            .O(N__22326),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    CascadeMux I__2172 (
            .O(N__22323),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ));
    InMux I__2171 (
            .O(N__22320),
            .I(N__22317));
    LocalMux I__2170 (
            .O(N__22317),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__2169 (
            .O(N__22314),
            .I(N__22311));
    LocalMux I__2168 (
            .O(N__22311),
            .I(N__22308));
    Odrv4 I__2167 (
            .O(N__22308),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    InMux I__2166 (
            .O(N__22305),
            .I(N__22302));
    LocalMux I__2165 (
            .O(N__22302),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ));
    InMux I__2164 (
            .O(N__22299),
            .I(N__22296));
    LocalMux I__2163 (
            .O(N__22296),
            .I(N__22293));
    Odrv4 I__2162 (
            .O(N__22293),
            .I(\current_shift_inst.PI_CTRL.N_46_21 ));
    InMux I__2161 (
            .O(N__22290),
            .I(N__22287));
    LocalMux I__2160 (
            .O(N__22287),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__2159 (
            .O(N__22284),
            .I(\current_shift_inst.control_input_cry_26 ));
    InMux I__2158 (
            .O(N__22281),
            .I(\current_shift_inst.control_input_cry_27 ));
    InMux I__2157 (
            .O(N__22278),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__2156 (
            .O(N__22275),
            .I(\current_shift_inst.control_input_cry_29 ));
    CascadeMux I__2155 (
            .O(N__22272),
            .I(\current_shift_inst.control_input_31_cascade_ ));
    InMux I__2154 (
            .O(N__22269),
            .I(N__22266));
    LocalMux I__2153 (
            .O(N__22266),
            .I(N__22263));
    Span4Mux_v I__2152 (
            .O(N__22263),
            .I(N__22260));
    Odrv4 I__2151 (
            .O(N__22260),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__2150 (
            .O(N__22257),
            .I(N__22254));
    LocalMux I__2149 (
            .O(N__22254),
            .I(N__22251));
    Odrv4 I__2148 (
            .O(N__22251),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ));
    CascadeMux I__2147 (
            .O(N__22248),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    CascadeMux I__2146 (
            .O(N__22245),
            .I(N__22240));
    InMux I__2145 (
            .O(N__22244),
            .I(N__22237));
    InMux I__2144 (
            .O(N__22243),
            .I(N__22234));
    InMux I__2143 (
            .O(N__22240),
            .I(N__22231));
    LocalMux I__2142 (
            .O(N__22237),
            .I(\current_shift_inst.N_1571_i ));
    LocalMux I__2141 (
            .O(N__22234),
            .I(\current_shift_inst.N_1571_i ));
    LocalMux I__2140 (
            .O(N__22231),
            .I(\current_shift_inst.N_1571_i ));
    InMux I__2139 (
            .O(N__22224),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__2138 (
            .O(N__22221),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__2137 (
            .O(N__22218),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__2136 (
            .O(N__22215),
            .I(\current_shift_inst.control_input_cry_20 ));
    InMux I__2135 (
            .O(N__22212),
            .I(\current_shift_inst.control_input_cry_21 ));
    InMux I__2134 (
            .O(N__22209),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__2133 (
            .O(N__22206),
            .I(bfn_3_14_0_));
    InMux I__2132 (
            .O(N__22203),
            .I(\current_shift_inst.control_input_cry_24 ));
    InMux I__2131 (
            .O(N__22200),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__2130 (
            .O(N__22197),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__2129 (
            .O(N__22194),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__2128 (
            .O(N__22191),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__2127 (
            .O(N__22188),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__2126 (
            .O(N__22185),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__2125 (
            .O(N__22182),
            .I(\current_shift_inst.control_input_cry_13 ));
    InMux I__2124 (
            .O(N__22179),
            .I(\current_shift_inst.control_input_cry_14 ));
    InMux I__2123 (
            .O(N__22176),
            .I(bfn_3_13_0_));
    InMux I__2122 (
            .O(N__22173),
            .I(\current_shift_inst.control_input_cry_16 ));
    InMux I__2121 (
            .O(N__22170),
            .I(N__22167));
    LocalMux I__2120 (
            .O(N__22167),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__2119 (
            .O(N__22164),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__2118 (
            .O(N__22161),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__2117 (
            .O(N__22158),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__2116 (
            .O(N__22155),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__2115 (
            .O(N__22152),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__2114 (
            .O(N__22149),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__2113 (
            .O(N__22146),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__2112 (
            .O(N__22143),
            .I(bfn_3_12_0_));
    InMux I__2111 (
            .O(N__22140),
            .I(N__22137));
    LocalMux I__2110 (
            .O(N__22137),
            .I(N__22134));
    Odrv12 I__2109 (
            .O(N__22134),
            .I(un8_start_stop));
    InMux I__2108 (
            .O(N__22131),
            .I(N__22128));
    LocalMux I__2107 (
            .O(N__22128),
            .I(N__22125));
    Odrv4 I__2106 (
            .O(N__22125),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    CascadeMux I__2105 (
            .O(N__22122),
            .I(N__22119));
    InMux I__2104 (
            .O(N__22119),
            .I(N__22116));
    LocalMux I__2103 (
            .O(N__22116),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__2102 (
            .O(N__22113),
            .I(N__22110));
    LocalMux I__2101 (
            .O(N__22110),
            .I(N__22107));
    Odrv4 I__2100 (
            .O(N__22107),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__2099 (
            .O(N__22104),
            .I(N__22101));
    LocalMux I__2098 (
            .O(N__22101),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__2097 (
            .O(N__22098),
            .I(N__22095));
    LocalMux I__2096 (
            .O(N__22095),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__2095 (
            .O(N__22092),
            .I(N__22089));
    LocalMux I__2094 (
            .O(N__22089),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__2093 (
            .O(N__22086),
            .I(N__22083));
    LocalMux I__2092 (
            .O(N__22083),
            .I(N__22080));
    Odrv4 I__2091 (
            .O(N__22080),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__2090 (
            .O(N__22077),
            .I(N__22074));
    LocalMux I__2089 (
            .O(N__22074),
            .I(N__22071));
    Odrv4 I__2088 (
            .O(N__22071),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    CascadeMux I__2087 (
            .O(N__22068),
            .I(N__22065));
    InMux I__2086 (
            .O(N__22065),
            .I(N__22062));
    LocalMux I__2085 (
            .O(N__22062),
            .I(N__22059));
    Span4Mux_v I__2084 (
            .O(N__22059),
            .I(N__22056));
    Odrv4 I__2083 (
            .O(N__22056),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__2082 (
            .O(N__22053),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__2081 (
            .O(N__22050),
            .I(N__22047));
    LocalMux I__2080 (
            .O(N__22047),
            .I(N__22044));
    Odrv4 I__2079 (
            .O(N__22044),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__2078 (
            .O(N__22041),
            .I(N__22038));
    LocalMux I__2077 (
            .O(N__22038),
            .I(N__22035));
    Odrv4 I__2076 (
            .O(N__22035),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__2075 (
            .O(N__22032),
            .I(N__22029));
    LocalMux I__2074 (
            .O(N__22029),
            .I(N__22026));
    Odrv4 I__2073 (
            .O(N__22026),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__2072 (
            .O(N__22023),
            .I(N__22020));
    LocalMux I__2071 (
            .O(N__22020),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__2070 (
            .O(N__22017),
            .I(N__22014));
    LocalMux I__2069 (
            .O(N__22014),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__2068 (
            .O(N__22011),
            .I(N__22008));
    LocalMux I__2067 (
            .O(N__22008),
            .I(N__22005));
    Odrv4 I__2066 (
            .O(N__22005),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__2065 (
            .O(N__22002),
            .I(N__21999));
    LocalMux I__2064 (
            .O(N__21999),
            .I(N__21996));
    Odrv4 I__2063 (
            .O(N__21996),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__2062 (
            .O(N__21993),
            .I(N__21990));
    LocalMux I__2061 (
            .O(N__21990),
            .I(N__21987));
    Glb2LocalMux I__2060 (
            .O(N__21987),
            .I(N__21984));
    GlobalMux I__2059 (
            .O(N__21984),
            .I(clk_12mhz));
    IoInMux I__2058 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__2057 (
            .O(N__21978),
            .I(N__21975));
    Span4Mux_s0_v I__2056 (
            .O(N__21975),
            .I(N__21972));
    Span4Mux_h I__2055 (
            .O(N__21972),
            .I(N__21969));
    Odrv4 I__2054 (
            .O(N__21969),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    CascadeMux I__2053 (
            .O(N__21966),
            .I(N__21963));
    InMux I__2052 (
            .O(N__21963),
            .I(N__21960));
    LocalMux I__2051 (
            .O(N__21960),
            .I(N__21957));
    Odrv4 I__2050 (
            .O(N__21957),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__2049 (
            .O(N__21954),
            .I(N__21951));
    LocalMux I__2048 (
            .O(N__21951),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__2047 (
            .O(N__21948),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__2046 (
            .O(N__21945),
            .I(N__21942));
    InMux I__2045 (
            .O(N__21942),
            .I(N__21939));
    LocalMux I__2044 (
            .O(N__21939),
            .I(N__21936));
    Odrv4 I__2043 (
            .O(N__21936),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__2042 (
            .O(N__21933),
            .I(N__21930));
    LocalMux I__2041 (
            .O(N__21930),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__2040 (
            .O(N__21927),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__2039 (
            .O(N__21924),
            .I(N__21921));
    InMux I__2038 (
            .O(N__21921),
            .I(N__21918));
    LocalMux I__2037 (
            .O(N__21918),
            .I(N__21915));
    Span4Mux_v I__2036 (
            .O(N__21915),
            .I(N__21912));
    Odrv4 I__2035 (
            .O(N__21912),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__2034 (
            .O(N__21909),
            .I(bfn_2_13_0_));
    CascadeMux I__2033 (
            .O(N__21906),
            .I(N__21903));
    InMux I__2032 (
            .O(N__21903),
            .I(N__21900));
    LocalMux I__2031 (
            .O(N__21900),
            .I(N__21897));
    Span4Mux_v I__2030 (
            .O(N__21897),
            .I(N__21894));
    Odrv4 I__2029 (
            .O(N__21894),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__2028 (
            .O(N__21891),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__2027 (
            .O(N__21888),
            .I(N__21885));
    InMux I__2026 (
            .O(N__21885),
            .I(N__21882));
    LocalMux I__2025 (
            .O(N__21882),
            .I(N__21879));
    Span4Mux_v I__2024 (
            .O(N__21879),
            .I(N__21876));
    Odrv4 I__2023 (
            .O(N__21876),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__2022 (
            .O(N__21873),
            .I(N__21870));
    LocalMux I__2021 (
            .O(N__21870),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__2020 (
            .O(N__21867),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__2019 (
            .O(N__21864),
            .I(N__21861));
    LocalMux I__2018 (
            .O(N__21861),
            .I(N__21858));
    Odrv4 I__2017 (
            .O(N__21858),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__2016 (
            .O(N__21855),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__2015 (
            .O(N__21852),
            .I(N__21849));
    InMux I__2014 (
            .O(N__21849),
            .I(N__21846));
    LocalMux I__2013 (
            .O(N__21846),
            .I(N__21843));
    Odrv4 I__2012 (
            .O(N__21843),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__2011 (
            .O(N__21840),
            .I(N__21837));
    LocalMux I__2010 (
            .O(N__21837),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__2009 (
            .O(N__21834),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__2008 (
            .O(N__21831),
            .I(N__21828));
    InMux I__2007 (
            .O(N__21828),
            .I(N__21825));
    LocalMux I__2006 (
            .O(N__21825),
            .I(N__21822));
    Span4Mux_v I__2005 (
            .O(N__21822),
            .I(N__21819));
    Odrv4 I__2004 (
            .O(N__21819),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__2003 (
            .O(N__21816),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    CascadeMux I__2002 (
            .O(N__21813),
            .I(N__21810));
    InMux I__2001 (
            .O(N__21810),
            .I(N__21807));
    LocalMux I__2000 (
            .O(N__21807),
            .I(N__21804));
    Span4Mux_v I__1999 (
            .O(N__21804),
            .I(N__21801));
    Odrv4 I__1998 (
            .O(N__21801),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1997 (
            .O(N__21798),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__1996 (
            .O(N__21795),
            .I(N__21792));
    InMux I__1995 (
            .O(N__21792),
            .I(N__21789));
    LocalMux I__1994 (
            .O(N__21789),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1993 (
            .O(N__21786),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__1992 (
            .O(N__21783),
            .I(N__21780));
    InMux I__1991 (
            .O(N__21780),
            .I(N__21777));
    LocalMux I__1990 (
            .O(N__21777),
            .I(N__21774));
    Span4Mux_v I__1989 (
            .O(N__21774),
            .I(N__21771));
    Odrv4 I__1988 (
            .O(N__21771),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__1987 (
            .O(N__21768),
            .I(N__21765));
    LocalMux I__1986 (
            .O(N__21765),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__1985 (
            .O(N__21762),
            .I(bfn_2_12_0_));
    CascadeMux I__1984 (
            .O(N__21759),
            .I(N__21756));
    InMux I__1983 (
            .O(N__21756),
            .I(N__21753));
    LocalMux I__1982 (
            .O(N__21753),
            .I(N__21750));
    Odrv4 I__1981 (
            .O(N__21750),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1980 (
            .O(N__21747),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1979 (
            .O(N__21744),
            .I(N__21741));
    InMux I__1978 (
            .O(N__21741),
            .I(N__21738));
    LocalMux I__1977 (
            .O(N__21738),
            .I(N__21735));
    Span4Mux_v I__1976 (
            .O(N__21735),
            .I(N__21732));
    Odrv4 I__1975 (
            .O(N__21732),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1974 (
            .O(N__21729),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__1973 (
            .O(N__21726),
            .I(N__21723));
    LocalMux I__1972 (
            .O(N__21723),
            .I(N__21720));
    Odrv4 I__1971 (
            .O(N__21720),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1970 (
            .O(N__21717),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1969 (
            .O(N__21714),
            .I(N__21711));
    InMux I__1968 (
            .O(N__21711),
            .I(N__21708));
    LocalMux I__1967 (
            .O(N__21708),
            .I(N__21705));
    Odrv4 I__1966 (
            .O(N__21705),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1965 (
            .O(N__21702),
            .I(N__21699));
    LocalMux I__1964 (
            .O(N__21699),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__1963 (
            .O(N__21696),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__1962 (
            .O(N__21693),
            .I(N__21690));
    InMux I__1961 (
            .O(N__21690),
            .I(N__21687));
    LocalMux I__1960 (
            .O(N__21687),
            .I(N__21684));
    Span4Mux_v I__1959 (
            .O(N__21684),
            .I(N__21681));
    Odrv4 I__1958 (
            .O(N__21681),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1957 (
            .O(N__21678),
            .I(N__21675));
    LocalMux I__1956 (
            .O(N__21675),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__1955 (
            .O(N__21672),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__1954 (
            .O(N__21669),
            .I(N__21666));
    InMux I__1953 (
            .O(N__21666),
            .I(N__21663));
    LocalMux I__1952 (
            .O(N__21663),
            .I(N__21660));
    Odrv4 I__1951 (
            .O(N__21660),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1950 (
            .O(N__21657),
            .I(N__21654));
    LocalMux I__1949 (
            .O(N__21654),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__1948 (
            .O(N__21651),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1947 (
            .O(N__21648),
            .I(N__21645));
    InMux I__1946 (
            .O(N__21645),
            .I(N__21642));
    LocalMux I__1945 (
            .O(N__21642),
            .I(N__21639));
    Span4Mux_h I__1944 (
            .O(N__21639),
            .I(N__21636));
    Odrv4 I__1943 (
            .O(N__21636),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1942 (
            .O(N__21633),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__1941 (
            .O(N__21630),
            .I(N__21627));
    InMux I__1940 (
            .O(N__21627),
            .I(N__21624));
    LocalMux I__1939 (
            .O(N__21624),
            .I(N__21621));
    Odrv4 I__1938 (
            .O(N__21621),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__1937 (
            .O(N__21618),
            .I(N__21615));
    LocalMux I__1936 (
            .O(N__21615),
            .I(N__21612));
    Odrv4 I__1935 (
            .O(N__21612),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__1934 (
            .O(N__21609),
            .I(bfn_2_11_0_));
    InMux I__1933 (
            .O(N__21606),
            .I(N__21603));
    LocalMux I__1932 (
            .O(N__21603),
            .I(N__21600));
    Odrv12 I__1931 (
            .O(N__21600),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1930 (
            .O(N__21597),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__1929 (
            .O(N__21594),
            .I(N__21591));
    InMux I__1928 (
            .O(N__21591),
            .I(N__21588));
    LocalMux I__1927 (
            .O(N__21588),
            .I(N__21585));
    Odrv4 I__1926 (
            .O(N__21585),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1925 (
            .O(N__21582),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__1924 (
            .O(N__21579),
            .I(N__21576));
    LocalMux I__1923 (
            .O(N__21576),
            .I(N__21573));
    Odrv4 I__1922 (
            .O(N__21573),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__1921 (
            .O(N__21570),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1920 (
            .O(N__21567),
            .I(N__21564));
    InMux I__1919 (
            .O(N__21564),
            .I(N__21561));
    LocalMux I__1918 (
            .O(N__21561),
            .I(N__21558));
    Odrv12 I__1917 (
            .O(N__21558),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1916 (
            .O(N__21555),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__1915 (
            .O(N__21552),
            .I(N__21549));
    InMux I__1914 (
            .O(N__21549),
            .I(N__21546));
    LocalMux I__1913 (
            .O(N__21546),
            .I(N__21543));
    Odrv12 I__1912 (
            .O(N__21543),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1911 (
            .O(N__21540),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    InMux I__1910 (
            .O(N__21537),
            .I(N__21534));
    LocalMux I__1909 (
            .O(N__21534),
            .I(N__21531));
    Span4Mux_h I__1908 (
            .O(N__21531),
            .I(N__21528));
    Odrv4 I__1907 (
            .O(N__21528),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    CascadeMux I__1906 (
            .O(N__21525),
            .I(N__21519));
    CascadeMux I__1905 (
            .O(N__21524),
            .I(N__21515));
    InMux I__1904 (
            .O(N__21523),
            .I(N__21512));
    InMux I__1903 (
            .O(N__21522),
            .I(N__21496));
    InMux I__1902 (
            .O(N__21519),
            .I(N__21496));
    InMux I__1901 (
            .O(N__21518),
            .I(N__21496));
    InMux I__1900 (
            .O(N__21515),
            .I(N__21496));
    LocalMux I__1899 (
            .O(N__21512),
            .I(N__21493));
    CascadeMux I__1898 (
            .O(N__21511),
            .I(N__21490));
    CascadeMux I__1897 (
            .O(N__21510),
            .I(N__21487));
    CascadeMux I__1896 (
            .O(N__21509),
            .I(N__21484));
    CascadeMux I__1895 (
            .O(N__21508),
            .I(N__21481));
    CascadeMux I__1894 (
            .O(N__21507),
            .I(N__21478));
    CascadeMux I__1893 (
            .O(N__21506),
            .I(N__21475));
    CascadeMux I__1892 (
            .O(N__21505),
            .I(N__21472));
    LocalMux I__1891 (
            .O(N__21496),
            .I(N__21469));
    Span4Mux_h I__1890 (
            .O(N__21493),
            .I(N__21466));
    InMux I__1889 (
            .O(N__21490),
            .I(N__21459));
    InMux I__1888 (
            .O(N__21487),
            .I(N__21459));
    InMux I__1887 (
            .O(N__21484),
            .I(N__21459));
    InMux I__1886 (
            .O(N__21481),
            .I(N__21450));
    InMux I__1885 (
            .O(N__21478),
            .I(N__21450));
    InMux I__1884 (
            .O(N__21475),
            .I(N__21450));
    InMux I__1883 (
            .O(N__21472),
            .I(N__21450));
    Span4Mux_v I__1882 (
            .O(N__21469),
            .I(N__21447));
    Odrv4 I__1881 (
            .O(N__21466),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1880 (
            .O(N__21459),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    LocalMux I__1879 (
            .O(N__21450),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    Odrv4 I__1878 (
            .O(N__21447),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    CascadeMux I__1877 (
            .O(N__21438),
            .I(N__21435));
    InMux I__1876 (
            .O(N__21435),
            .I(N__21432));
    LocalMux I__1875 (
            .O(N__21432),
            .I(N__21429));
    Odrv4 I__1874 (
            .O(N__21429),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__1873 (
            .O(N__21426),
            .I(N__21423));
    InMux I__1872 (
            .O(N__21423),
            .I(N__21420));
    LocalMux I__1871 (
            .O(N__21420),
            .I(N__21417));
    Odrv12 I__1870 (
            .O(N__21417),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1869 (
            .O(N__21414),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__1868 (
            .O(N__21411),
            .I(N__21408));
    InMux I__1867 (
            .O(N__21408),
            .I(N__21405));
    LocalMux I__1866 (
            .O(N__21405),
            .I(N__21402));
    Odrv12 I__1865 (
            .O(N__21402),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1864 (
            .O(N__21399),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__1863 (
            .O(N__21396),
            .I(N__21393));
    InMux I__1862 (
            .O(N__21393),
            .I(N__21390));
    LocalMux I__1861 (
            .O(N__21390),
            .I(N__21387));
    Odrv4 I__1860 (
            .O(N__21387),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__1859 (
            .O(N__21384),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__1858 (
            .O(N__21381),
            .I(N__21378));
    InMux I__1857 (
            .O(N__21378),
            .I(N__21375));
    LocalMux I__1856 (
            .O(N__21375),
            .I(N__21372));
    Odrv12 I__1855 (
            .O(N__21372),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1854 (
            .O(N__21369),
            .I(N__21366));
    LocalMux I__1853 (
            .O(N__21366),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__1852 (
            .O(N__21363),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__1851 (
            .O(N__21360),
            .I(N__21357));
    InMux I__1850 (
            .O(N__21357),
            .I(N__21354));
    LocalMux I__1849 (
            .O(N__21354),
            .I(N__21351));
    Span4Mux_h I__1848 (
            .O(N__21351),
            .I(N__21348));
    Odrv4 I__1847 (
            .O(N__21348),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1846 (
            .O(N__21345),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    InMux I__1845 (
            .O(N__21342),
            .I(N__21339));
    LocalMux I__1844 (
            .O(N__21339),
            .I(N__21336));
    Span4Mux_v I__1843 (
            .O(N__21336),
            .I(N__21333));
    Odrv4 I__1842 (
            .O(N__21333),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__1841 (
            .O(N__21330),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1840 (
            .O(N__21327),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__1839 (
            .O(N__21324),
            .I(N__21321));
    LocalMux I__1838 (
            .O(N__21321),
            .I(N_94_i_i));
    InMux I__1837 (
            .O(N__21318),
            .I(N__21315));
    LocalMux I__1836 (
            .O(N__21315),
            .I(N__21312));
    Span4Mux_v I__1835 (
            .O(N__21312),
            .I(N__21309));
    Odrv4 I__1834 (
            .O(N__21309),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1833 (
            .O(N__21306),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    CascadeMux I__1832 (
            .O(N__21303),
            .I(N__21300));
    InMux I__1831 (
            .O(N__21300),
            .I(N__21297));
    LocalMux I__1830 (
            .O(N__21297),
            .I(N__21294));
    Span4Mux_v I__1829 (
            .O(N__21294),
            .I(N__21291));
    Odrv4 I__1828 (
            .O(N__21291),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1827 (
            .O(N__21288),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__1826 (
            .O(N__21285),
            .I(N__21282));
    LocalMux I__1825 (
            .O(N__21282),
            .I(N__21279));
    Span4Mux_v I__1824 (
            .O(N__21279),
            .I(N__21276));
    Odrv4 I__1823 (
            .O(N__21276),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1822 (
            .O(N__21273),
            .I(bfn_1_11_0_));
    InMux I__1821 (
            .O(N__21270),
            .I(N__21267));
    LocalMux I__1820 (
            .O(N__21267),
            .I(N__21264));
    Span4Mux_v I__1819 (
            .O(N__21264),
            .I(N__21261));
    Odrv4 I__1818 (
            .O(N__21261),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1817 (
            .O(N__21258),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1816 (
            .O(N__21255),
            .I(N__21252));
    LocalMux I__1815 (
            .O(N__21252),
            .I(N__21249));
    Span4Mux_v I__1814 (
            .O(N__21249),
            .I(N__21246));
    Odrv4 I__1813 (
            .O(N__21246),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1812 (
            .O(N__21243),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1811 (
            .O(N__21240),
            .I(N__21237));
    LocalMux I__1810 (
            .O(N__21237),
            .I(N__21234));
    Span4Mux_v I__1809 (
            .O(N__21234),
            .I(N__21231));
    Odrv4 I__1808 (
            .O(N__21231),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1807 (
            .O(N__21228),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1806 (
            .O(N__21225),
            .I(N__21222));
    LocalMux I__1805 (
            .O(N__21222),
            .I(N__21219));
    Span4Mux_v I__1804 (
            .O(N__21219),
            .I(N__21216));
    Odrv4 I__1803 (
            .O(N__21216),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1802 (
            .O(N__21213),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1801 (
            .O(N__21210),
            .I(N__21207));
    LocalMux I__1800 (
            .O(N__21207),
            .I(N__21204));
    Span4Mux_v I__1799 (
            .O(N__21204),
            .I(N__21201));
    Odrv4 I__1798 (
            .O(N__21201),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1797 (
            .O(N__21198),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1796 (
            .O(N__21195),
            .I(N__21192));
    LocalMux I__1795 (
            .O(N__21192),
            .I(N__21189));
    Span4Mux_v I__1794 (
            .O(N__21189),
            .I(N__21186));
    Odrv4 I__1793 (
            .O(N__21186),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1792 (
            .O(N__21183),
            .I(N__21180));
    InMux I__1791 (
            .O(N__21180),
            .I(N__21177));
    LocalMux I__1790 (
            .O(N__21177),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__1789 (
            .O(N__21174),
            .I(N__21171));
    LocalMux I__1788 (
            .O(N__21171),
            .I(N__21168));
    Span4Mux_v I__1787 (
            .O(N__21168),
            .I(N__21165));
    Odrv4 I__1786 (
            .O(N__21165),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1785 (
            .O(N__21162),
            .I(N__21159));
    InMux I__1784 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__1783 (
            .O(N__21156),
            .I(N__21153));
    Odrv4 I__1782 (
            .O(N__21153),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1781 (
            .O(N__21150),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1780 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__1779 (
            .O(N__21144),
            .I(N__21141));
    Span4Mux_v I__1778 (
            .O(N__21141),
            .I(N__21138));
    Odrv4 I__1777 (
            .O(N__21138),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1776 (
            .O(N__21135),
            .I(N__21132));
    InMux I__1775 (
            .O(N__21132),
            .I(N__21129));
    LocalMux I__1774 (
            .O(N__21129),
            .I(N__21126));
    Odrv4 I__1773 (
            .O(N__21126),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1772 (
            .O(N__21123),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__1771 (
            .O(N__21120),
            .I(N__21117));
    LocalMux I__1770 (
            .O(N__21117),
            .I(N__21114));
    Span4Mux_v I__1769 (
            .O(N__21114),
            .I(N__21111));
    Odrv4 I__1768 (
            .O(N__21111),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1767 (
            .O(N__21108),
            .I(N__21105));
    InMux I__1766 (
            .O(N__21105),
            .I(N__21102));
    LocalMux I__1765 (
            .O(N__21102),
            .I(N__21099));
    Odrv4 I__1764 (
            .O(N__21099),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1763 (
            .O(N__21096),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__1762 (
            .O(N__21093),
            .I(N__21090));
    LocalMux I__1761 (
            .O(N__21090),
            .I(N__21087));
    Span4Mux_v I__1760 (
            .O(N__21087),
            .I(N__21084));
    Odrv4 I__1759 (
            .O(N__21084),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1758 (
            .O(N__21081),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    CascadeMux I__1757 (
            .O(N__21078),
            .I(N__21075));
    InMux I__1756 (
            .O(N__21075),
            .I(N__21072));
    LocalMux I__1755 (
            .O(N__21072),
            .I(N__21069));
    Span4Mux_v I__1754 (
            .O(N__21069),
            .I(N__21066));
    Odrv4 I__1753 (
            .O(N__21066),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1752 (
            .O(N__21063),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    IoInMux I__1751 (
            .O(N__21060),
            .I(N__21057));
    LocalMux I__1750 (
            .O(N__21057),
            .I(N__21054));
    Span4Mux_s3_v I__1749 (
            .O(N__21054),
            .I(N__21051));
    Span4Mux_h I__1748 (
            .O(N__21051),
            .I(N__21048));
    Sp12to4 I__1747 (
            .O(N__21048),
            .I(N__21045));
    Span12Mux_v I__1746 (
            .O(N__21045),
            .I(N__21042));
    Span12Mux_v I__1745 (
            .O(N__21042),
            .I(N__21039));
    Odrv12 I__1744 (
            .O(N__21039),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1743 (
            .O(N__21036),
            .I(N__21033));
    LocalMux I__1742 (
            .O(N__21033),
            .I(N__21030));
    IoSpan4Mux I__1741 (
            .O(N__21030),
            .I(N__21027));
    IoSpan4Mux I__1740 (
            .O(N__21027),
            .I(N__21024));
    Odrv4 I__1739 (
            .O(N__21024),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_28_0_));
    defparam IN_MUX_bfv_15_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_29_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_15_29_0_));
    defparam IN_MUX_bfv_15_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_30_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_15_30_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_16_28_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_28_0_));
    defparam IN_MUX_bfv_16_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_29_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_16_29_0_));
    defparam IN_MUX_bfv_16_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_30_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_16_30_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_17_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_27_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_0_cry_7 ),
            .carryinitout(bfn_17_27_0_));
    defparam IN_MUX_bfv_20_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_25_0_));
    defparam IN_MUX_bfv_20_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_26_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_20_26_0_));
    defparam IN_MUX_bfv_20_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_27_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_20_27_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_30 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_7 ),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_15 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_23 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_30 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_7 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_15 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_23 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_11_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_25_0_));
    defparam IN_MUX_bfv_11_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .carryinitout(bfn_11_26_0_));
    defparam IN_MUX_bfv_11_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_27_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .carryinitout(bfn_11_27_0_));
    defparam IN_MUX_bfv_11_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_28_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_30 ),
            .carryinitout(bfn_11_28_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_12_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_27_0_));
    defparam IN_MUX_bfv_12_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_28_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_7 ),
            .carryinitout(bfn_12_28_0_));
    defparam IN_MUX_bfv_12_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_29_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_15 ),
            .carryinitout(bfn_12_29_0_));
    defparam IN_MUX_bfv_12_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_30_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_23 ),
            .carryinitout(bfn_12_30_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_30 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_7 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_15 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_23 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_5_14_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21060),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21036),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \phase_controller_inst1.stoper_tr.running_RNI6D081_0  (
            .USERSIGNALTOGLOBALBUFFER(N__31470),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst1.stoper_tr.un2_start_0_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.running_RNI96ON_0  (
            .USERSIGNALTOGLOBALBUFFER(N__28083),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un2_start_0_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__38226),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_153_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__46576),
            .CLKHFEN(N__46578),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__46577),
            .RGB2PWM(N__21324),
            .RGB1(rgb_g),
            .CURREN(N__46828),
            .RGB2(rgb_b),
            .RGB1PWM(N__22140),
            .RGB0PWM(N__52089),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_6_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_6_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_6_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_1_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_1_9_2 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_1_9_2  (
            .in0(N__31641),
            .in1(N__21369),
            .in2(_gnd_net_),
            .in3(N__22597),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52500),
            .ce(),
            .sr(N__51989));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_1_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_1_9_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_1_9_5  (
            .in0(N__22596),
            .in1(N__21618),
            .in2(_gnd_net_),
            .in3(N__31642),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52500),
            .ce(),
            .sr(N__51989));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__21195),
            .in2(N__21183),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__21174),
            .in2(N__21162),
            .in3(N__21150),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__21147),
            .in2(N__21135),
            .in3(N__21123),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__21120),
            .in2(N__21108),
            .in3(N__21096),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__21093),
            .in2(N__21524),
            .in3(N__21081),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__21518),
            .in2(N__21078),
            .in3(N__21063),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__21318),
            .in2(N__21525),
            .in3(N__21306),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__21522),
            .in2(N__21303),
            .in3(N__21288),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__21285),
            .in2(N__21505),
            .in3(N__21273),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__21270),
            .in2(N__21509),
            .in3(N__21258),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__21255),
            .in2(N__21506),
            .in3(N__21243),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__21240),
            .in2(N__21510),
            .in3(N__21228),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__21225),
            .in2(N__21507),
            .in3(N__21213),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__21210),
            .in2(N__21511),
            .in3(N__21198),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__21342),
            .in2(N__21508),
            .in3(N__21330),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21327),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_1_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_1_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_1_12_2  (
            .in0(N__22621),
            .in1(N__31589),
            .in2(_gnd_net_),
            .in3(N__21768),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52494),
            .ce(),
            .sr(N__52007));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_1_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_1_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_1_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_1_12_6  (
            .in0(N__22622),
            .in1(N__31590),
            .in2(_gnd_net_),
            .in3(N__21678),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52494),
            .ce(),
            .sr(N__52007));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_1_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_1_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_1_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_1_12_7  (
            .in0(N__31588),
            .in1(N__22623),
            .in2(_gnd_net_),
            .in3(N__21954),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52494),
            .ce(),
            .sr(N__52007));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_1_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_1_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_1_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_1_13_1  (
            .in0(N__22624),
            .in1(N__31592),
            .in2(_gnd_net_),
            .in3(N__21702),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52491),
            .ce(),
            .sr(N__52014));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_1_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_1_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_1_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_1_13_3  (
            .in0(N__22625),
            .in1(N__31593),
            .in2(_gnd_net_),
            .in3(N__21933),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52491),
            .ce(),
            .sr(N__52014));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_1_13_5  (
            .in0(N__22626),
            .in1(N__31594),
            .in2(_gnd_net_),
            .in3(N__21873),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52491),
            .ce(),
            .sr(N__52014));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_14_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_1_14_5  (
            .in0(N__31591),
            .in1(N__22646),
            .in2(_gnd_net_),
            .in3(N__21840),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52485),
            .ce(),
            .sr(N__52023));
    defparam \phase_controller_inst1.N_94_i_i_LC_1_30_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_94_i_i_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_94_i_i_LC_1_30_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_94_i_i_LC_1_30_2  (
            .in0(N__52088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36612),
            .lcout(N_94_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_2_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_2_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__21537),
            .in2(_gnd_net_),
            .in3(N__21523),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_2_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_2_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_2_9_1  (
            .in0(N__30232),
            .in1(N__30106),
            .in2(N__30928),
            .in3(N__30173),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_2_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_2_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_2_9_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_2_9_5  (
            .in0(N__31643),
            .in1(N__21657),
            .in2(_gnd_net_),
            .in3(N__22595),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52499),
            .ce(),
            .sr(N__51980));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_10_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__36681),
            .in2(N__21438),
            .in3(N__22628),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(N__52497),
            .ce(),
            .sr(N__51991));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_2_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_2_10_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_2_10_1  (
            .in0(N__22627),
            .in1(N__30427),
            .in2(N__21426),
            .in3(N__21414),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(N__52497),
            .ce(),
            .sr(N__51991));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_10_2 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_2_10_2  (
            .in0(N__22647),
            .in1(N__30351),
            .in2(N__21411),
            .in3(N__21399),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(N__52497),
            .ce(),
            .sr(N__51991));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__30295),
            .in2(N__21396),
            .in3(N__21384),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__30228),
            .in2(N__21381),
            .in3(N__21363),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__30171),
            .in2(N__21360),
            .in3(N__21345),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__30105),
            .in2(N__21669),
            .in3(N__21651),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__30057),
            .in2(N__21648),
            .in3(N__21633),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__30927),
            .in2(N__21630),
            .in3(N__21609),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__21606),
            .in2(N__30860),
            .in3(N__21597),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__30793),
            .in2(N__21594),
            .in3(N__21582),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__21579),
            .in2(N__30731),
            .in3(N__21570),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__30655),
            .in2(N__21567),
            .in3(N__21555),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__30598),
            .in2(N__21552),
            .in3(N__21540),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__30547),
            .in2(N__21813),
            .in3(N__21798),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__30478),
            .in2(N__21795),
            .in3(N__21786),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__31419),
            .in2(N__21783),
            .in3(N__21762),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__31360),
            .in2(N__21759),
            .in3(N__21747),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__31296),
            .in2(N__21744),
            .in3(N__21729),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__21726),
            .in2(N__31229),
            .in3(N__21717),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__31155),
            .in2(N__21714),
            .in3(N__21696),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__31101),
            .in2(N__21693),
            .in3(N__21672),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__31041),
            .in2(N__21966),
            .in3(N__21948),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__30981),
            .in2(N__21945),
            .in3(N__21927),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__32016),
            .in2(N__21924),
            .in3(N__21909),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__31954),
            .in2(N__21906),
            .in3(N__21891),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__31878),
            .in2(N__21888),
            .in3(N__21867),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__21864),
            .in2(N__31824),
            .in3(N__21855),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__31747),
            .in2(N__21852),
            .in3(N__21834),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__31689),
            .in2(N__21831),
            .in3(N__21816),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_2_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_2_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_er_31_LC_2_13_6  (
            .in0(N__22077),
            .in1(N__31595),
            .in2(N__22068),
            .in3(N__22053),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52486),
            .ce(N__22649),
            .sr(N__52008));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_0  (
            .in0(N__31582),
            .in1(N__22632),
            .in2(_gnd_net_),
            .in3(N__22050),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52482),
            .ce(),
            .sr(N__52015));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_14_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_2_14_1  (
            .in0(N__22041),
            .in1(N__31587),
            .in2(N__22652),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52482),
            .ce(),
            .sr(N__52015));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_2_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_2_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_2_14_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_2_14_3  (
            .in0(N__22032),
            .in1(_gnd_net_),
            .in2(N__22653),
            .in3(N__31584),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52482),
            .ce(),
            .sr(N__52015));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_2_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_2_14_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_2_14_4  (
            .in0(N__31583),
            .in1(N__22633),
            .in2(_gnd_net_),
            .in3(N__22023),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52482),
            .ce(),
            .sr(N__52015));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_2_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_2_14_5 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_2_14_5  (
            .in0(N__22017),
            .in1(N__31586),
            .in2(N__22651),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52482),
            .ce(),
            .sr(N__52015));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_7  (
            .in0(N__22011),
            .in1(N__31585),
            .in2(N__22650),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52482),
            .ce(),
            .sr(N__52015));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1  (
            .in0(N__31613),
            .in1(N__22002),
            .in2(_gnd_net_),
            .in3(N__22648),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52478),
            .ce(),
            .sr(N__52024));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_1.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21993),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un8_start_stop_LC_2_30_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.un8_start_stop_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un8_start_stop_LC_2_30_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.un8_start_stop_LC_2_30_2  (
            .in0(N__52087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36611),
            .lcout(un8_start_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_3_9_0  (
            .in0(N__22550),
            .in1(N__31650),
            .in2(_gnd_net_),
            .in3(N__22131),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52498),
            .ce(),
            .sr(N__51976));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_9_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_3_9_3  (
            .in0(N__31648),
            .in1(_gnd_net_),
            .in2(N__22122),
            .in3(N__22552),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52498),
            .ce(),
            .sr(N__51976));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_3_9_5  (
            .in0(N__31647),
            .in1(N__22113),
            .in2(_gnd_net_),
            .in3(N__22551),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52498),
            .ce(),
            .sr(N__51976));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_9_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_3_9_7  (
            .in0(N__31649),
            .in1(N__22104),
            .in2(_gnd_net_),
            .in3(N__22553),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52498),
            .ce(),
            .sr(N__51976));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_3_10_0  (
            .in0(N__22554),
            .in1(N__31652),
            .in2(_gnd_net_),
            .in3(N__22098),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52495),
            .ce(),
            .sr(N__51981));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_3_10_1  (
            .in0(N__31651),
            .in1(N__22092),
            .in2(_gnd_net_),
            .in3(N__22557),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52495),
            .ce(),
            .sr(N__51981));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_3_10_2  (
            .in0(N__22555),
            .in1(N__31653),
            .in2(_gnd_net_),
            .in3(N__22086),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52495),
            .ce(),
            .sr(N__51981));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_3_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_3_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_3_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(N__22244),
            .in2(_gnd_net_),
            .in3(N__23673),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52495),
            .ce(),
            .sr(N__51981));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_10_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_3_10_6  (
            .in0(N__22556),
            .in1(N__31654),
            .in2(_gnd_net_),
            .in3(N__22170),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52495),
            .ce(),
            .sr(N__51981));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_3_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_3_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__23669),
            .in2(N__22245),
            .in3(N__22243),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_3_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_3_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__23688),
            .in2(_gnd_net_),
            .in3(N__22164),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_3_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_3_11_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__22359),
            .in2(_gnd_net_),
            .in3(N__22161),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_3_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_3_11_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__23649),
            .in2(_gnd_net_),
            .in3(N__22158),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_3_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_3_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__23634),
            .in2(_gnd_net_),
            .in3(N__22155),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_3_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_3_11_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(N__22365),
            .in2(_gnd_net_),
            .in3(N__22152),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_3_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_3_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(N__22395),
            .in2(_gnd_net_),
            .in3(N__22149),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_3_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_3_11_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_3_11_7  (
            .in0(_gnd_net_),
            .in1(N__22371),
            .in2(_gnd_net_),
            .in3(N__22146),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_3_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_3_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__22377),
            .in2(_gnd_net_),
            .in3(N__22143),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_3_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_3_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(N__23586),
            .in2(_gnd_net_),
            .in3(N__22197),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_3_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_3_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(N__22455),
            .in2(_gnd_net_),
            .in3(N__22194),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_3_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_3_12_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(N__23598),
            .in2(_gnd_net_),
            .in3(N__22191),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_3_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_3_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(N__22353),
            .in2(_gnd_net_),
            .in3(N__22188),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_3_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_3_12_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_3_12_5  (
            .in0(_gnd_net_),
            .in1(N__22449),
            .in2(_gnd_net_),
            .in3(N__22185),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_3_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_3_12_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(N__23574),
            .in2(_gnd_net_),
            .in3(N__22182),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_3_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_3_12_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_3_12_7  (
            .in0(_gnd_net_),
            .in1(N__23529),
            .in2(_gnd_net_),
            .in3(N__22179),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_3_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_3_13_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__23700),
            .in2(_gnd_net_),
            .in3(N__22176),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_3_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_3_13_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__23541),
            .in2(_gnd_net_),
            .in3(N__22173),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_3_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_3_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(N__22443),
            .in2(_gnd_net_),
            .in3(N__22224),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_3_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_3_13_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(N__23931),
            .in2(_gnd_net_),
            .in3(N__22221),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_3_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_3_13_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__22437),
            .in2(_gnd_net_),
            .in3(N__22218),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_3_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_3_13_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(N__23553),
            .in2(_gnd_net_),
            .in3(N__22215),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_3_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_3_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(N__22407),
            .in2(_gnd_net_),
            .in3(N__22212),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_3_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_3_13_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__22719),
            .in2(_gnd_net_),
            .in3(N__22209),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_3_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_3_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__22401),
            .in2(_gnd_net_),
            .in3(N__22206),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_3_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_3_14_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__22713),
            .in2(_gnd_net_),
            .in3(N__22203),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_3_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_3_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__23562),
            .in2(_gnd_net_),
            .in3(N__22200),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_3_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_3_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__22413),
            .in2(_gnd_net_),
            .in3(N__22284),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_3_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_3_14_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__24414),
            .in2(_gnd_net_),
            .in3(N__22281),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_3_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_3_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__22695),
            .in2(_gnd_net_),
            .in3(N__22278),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_3_14_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_3_14_6  (
            .in0(N__24586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22275),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(\current_shift_inst.control_input_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_3_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_3_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22272),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_3_15_7  (
            .in0(N__31635),
            .in1(N__22269),
            .in2(_gnd_net_),
            .in3(N__22620),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52470),
            .ce(),
            .sr(N__52016));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_9_0 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_9_0  (
            .in0(N__30059),
            .in1(N__30296),
            .in2(N__30368),
            .in3(N__22257),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_4_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_4_9_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_4_9_1  (
            .in0(N__22686),
            .in1(N__22299),
            .in2(N__22248),
            .in3(N__22314),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_4_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_4_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24560),
            .lcout(\current_shift_inst.N_1571_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_10_3  (
            .in0(N__30597),
            .in1(N__30651),
            .in2(N__30794),
            .in3(N__30462),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_4_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_4_10_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_4_10_4  (
            .in0(N__30113),
            .in1(N__30172),
            .in2(_gnd_net_),
            .in3(N__30239),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_4_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_4_10_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_4_10_5  (
            .in0(N__30058),
            .in1(N__30929),
            .in2(N__22335),
            .in3(N__22332),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_10_7 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_10_7  (
            .in0(N__30352),
            .in1(N__30431),
            .in2(N__36697),
            .in3(N__30294),
            .lcout(\current_shift_inst.PI_CTRL.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_4_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_4_11_0  (
            .in0(N__30853),
            .in1(N__22389),
            .in2(N__30548),
            .in3(N__22290),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_4_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_4_11_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_4_11_1  (
            .in0(N__31636),
            .in1(N__31350),
            .in2(N__22326),
            .in3(N__22461),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_4_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_4_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_4_11_2  (
            .in0(N__22707),
            .in1(N__22422),
            .in2(N__22323),
            .in3(N__22320),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_4_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_4_11_4  (
            .in0(N__22431),
            .in1(N__22383),
            .in2(N__22347),
            .in3(N__22305),
            .lcout(\current_shift_inst.PI_CTRL.N_46_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_4_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_4_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_4_11_7  (
            .in0(N__31227),
            .in1(N__31429),
            .in2(N__31307),
            .in3(N__31114),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_4_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_4_12_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_4_12_0  (
            .in0(N__24639),
            .in1(N__24135),
            .in2(_gnd_net_),
            .in3(N__24563),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_4_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_4_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__31756),
            .in2(_gnd_net_),
            .in3(N__31042),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_4_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_4_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_4_12_2  (
            .in0(N__31757),
            .in1(N__30540),
            .in2(N__31049),
            .in3(N__30852),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_4_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_4_12_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_4_12_3  (
            .in0(N__24565),
            .in1(N__24858),
            .in2(_gnd_net_),
            .in3(N__24111),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_4_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_4_12_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_4_12_4  (
            .in0(N__24615),
            .in1(N__24123),
            .in2(_gnd_net_),
            .in3(N__24564),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_4_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_4_12_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_4_12_5  (
            .in0(N__24562),
            .in1(N__24147),
            .in2(_gnd_net_),
            .in3(N__24654),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_4_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_4_12_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_4_12_6  (
            .in0(N__24003),
            .in1(N__24693),
            .in2(_gnd_net_),
            .in3(N__24561),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_4_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_4_12_7 .LUT_INIT=16'b0000010111110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_4_12_7  (
            .in0(N__24792),
            .in1(_gnd_net_),
            .in2(N__24587),
            .in3(N__24267),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_4_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_4_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_4_13_0  (
            .in0(N__31825),
            .in1(N__31882),
            .in2(N__31706),
            .in3(N__30727),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_4_13_1 .LUT_INIT=16'b0001101100011011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_4_13_1  (
            .in0(N__24588),
            .in1(N__24825),
            .in2(N__24090),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_4_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_4_13_3 .LUT_INIT=16'b0011010100110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_4_13_3  (
            .in0(N__24774),
            .in1(N__24252),
            .in2(N__24594),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_4_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_4_13_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_4_13_4  (
            .in0(N__24592),
            .in1(N__24192),
            .in2(_gnd_net_),
            .in3(N__24996),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_4_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_4_13_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_4_13_5  (
            .in0(N__24963),
            .in1(N__24381),
            .in2(_gnd_net_),
            .in3(N__24593),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_4_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_4_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_4_13_6  (
            .in0(N__31156),
            .in1(N__32017),
            .in2(N__31958),
            .in3(N__30982),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_4_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_4_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_4_13_7  (
            .in0(N__32018),
            .in1(N__31953),
            .in2(N__30989),
            .in3(N__31157),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_4_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_4_14_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_4_14_0  (
            .in0(N__24288),
            .in1(N__24585),
            .in2(_gnd_net_),
            .in3(N__25098),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_4_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_4_14_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_4_14_2  (
            .in0(N__24348),
            .in1(N__24921),
            .in2(_gnd_net_),
            .in3(N__24581),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_4_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_4_14_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_4_14_3  (
            .in0(N__24583),
            .in1(N__24882),
            .in2(_gnd_net_),
            .in3(N__24324),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_4_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_4_14_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_4_14_5  (
            .in0(N__24582),
            .in1(N__24336),
            .in2(_gnd_net_),
            .in3(N__24903),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_4_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_4_14_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_4_14_6  (
            .in0(N__25146),
            .in1(N__24309),
            .in2(_gnd_net_),
            .in3(N__24584),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_4_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_4_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_4_14_7  (
            .in0(N__31690),
            .in1(N__31886),
            .in2(N__31826),
            .in3(N__30723),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_4_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_4_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24559),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_4_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_4_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_4_15_4  (
            .in0(N__31228),
            .in1(N__31303),
            .in2(N__31436),
            .in3(N__31115),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_46_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_4_15_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__31640),
            .in2(N__22689),
            .in3(N__31361),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22677),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52449),
            .ce(),
            .sr(N__52031));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4  (
            .in0(N__31655),
            .in1(N__22558),
            .in2(_gnd_net_),
            .in3(N__22473),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52492),
            .ce(),
            .sr(N__51970));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_10_4  (
            .in0(N__30602),
            .in1(N__30656),
            .in2(N__30482),
            .in3(N__30774),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__22824),
            .in2(_gnd_net_),
            .in3(N__22833),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_5_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_5_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__22818),
            .in2(_gnd_net_),
            .in3(N__22809),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_5_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_5_11_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22806),
            .in3(N__22794),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_5_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_5_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__22791),
            .in2(_gnd_net_),
            .in3(N__22782),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_5_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_5_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__22779),
            .in2(_gnd_net_),
            .in3(N__22770),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_5_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_5_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__22767),
            .in2(_gnd_net_),
            .in3(N__22758),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_5_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_5_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__22755),
            .in2(_gnd_net_),
            .in3(N__22746),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_5_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_5_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__22743),
            .in2(_gnd_net_),
            .in3(N__22734),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__52483),
            .ce(),
            .sr(N__51977));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_5_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_5_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__22731),
            .in2(_gnd_net_),
            .in3(N__22722),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_5_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_5_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__22932),
            .in2(_gnd_net_),
            .in3(N__22923),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_5_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_5_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__22920),
            .in2(_gnd_net_),
            .in3(N__22911),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_5_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_5_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22908),
            .in3(N__22896),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_5_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_5_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__22893),
            .in2(_gnd_net_),
            .in3(N__22884),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_5_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_5_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__22881),
            .in2(_gnd_net_),
            .in3(N__22872),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_5_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_5_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__22869),
            .in2(_gnd_net_),
            .in3(N__22860),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_5_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_5_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__22857),
            .in2(_gnd_net_),
            .in3(N__22848),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__52479),
            .ce(),
            .sr(N__51982));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_5_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_5_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__22845),
            .in2(_gnd_net_),
            .in3(N__22836),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_5_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_5_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__23040),
            .in2(_gnd_net_),
            .in3(N__23031),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_5_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_5_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__23028),
            .in2(_gnd_net_),
            .in3(N__23019),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_5_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_5_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__23016),
            .in2(_gnd_net_),
            .in3(N__23007),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_5_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_5_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__23004),
            .in2(_gnd_net_),
            .in3(N__22995),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_5_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_5_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__22992),
            .in2(_gnd_net_),
            .in3(N__22983),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_5_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_5_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__22980),
            .in2(_gnd_net_),
            .in3(N__22971),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_5_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_5_13_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22968),
            .in3(N__22956),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__52471),
            .ce(),
            .sr(N__51992));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_5_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_5_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__22953),
            .in2(_gnd_net_),
            .in3(N__22944),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_5_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_5_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__22941),
            .in2(_gnd_net_),
            .in3(N__23163),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_5_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_5_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__23160),
            .in2(_gnd_net_),
            .in3(N__23151),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_5_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_5_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__23148),
            .in2(_gnd_net_),
            .in3(N__23139),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_5_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_5_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__23136),
            .in2(_gnd_net_),
            .in3(N__23127),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_5_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_5_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__23124),
            .in2(_gnd_net_),
            .in3(N__23115),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_5_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_5_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__23112),
            .in2(_gnd_net_),
            .in3(N__23103),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_5_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__23100),
            .in2(_gnd_net_),
            .in3(N__23091),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52465),
            .ce(),
            .sr(N__51995));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23087),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52459),
            .ce(),
            .sr(N__52001));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23060),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52459),
            .ce(),
            .sr(N__52001));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_5_15_3  (
            .in0(N__23318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52459),
            .ce(),
            .sr(N__52001));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23298),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52455),
            .ce(),
            .sr(N__52009));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23279),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52455),
            .ce(),
            .sr(N__52009));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23255),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52455),
            .ce(),
            .sr(N__52009));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23231),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52455),
            .ce(),
            .sr(N__52009));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23207),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52450),
            .ce(),
            .sr(N__52017));
    defparam \phase_controller_inst1.start_flag_LC_5_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_flag_LC_5_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_flag_LC_5_17_2 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \phase_controller_inst1.start_flag_LC_5_17_2  (
            .in0(N__36588),
            .in1(N__36529),
            .in2(N__36512),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52450),
            .ce(),
            .sr(N__52017));
    defparam \phase_controller_inst1.state_4_LC_5_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_5_17_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_5_17_5 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \phase_controller_inst1.state_4_LC_5_17_5  (
            .in0(N__36530),
            .in1(N__36589),
            .in2(_gnd_net_),
            .in3(N__36505),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52450),
            .ce(),
            .sr(N__52017));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23183),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52450),
            .ce(),
            .sr(N__52017));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23516),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52442),
            .ce(),
            .sr(N__52025));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23489),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52442),
            .ce(),
            .sr(N__52025));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23459),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52436),
            .ce(),
            .sr(N__52032));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23435),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52436),
            .ce(),
            .sr(N__52032));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_5_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_5_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_5_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_5_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23415),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52431),
            .ce(),
            .sr(N__52036));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_5_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_5_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_5_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_5_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23399),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52425),
            .ce(),
            .sr(N__52041));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_5_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23378),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52425),
            .ce(),
            .sr(N__52041));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23354),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52420),
            .ce(),
            .sr(N__52044));
    defparam \delay_measurement_inst.start_timer_hc_LC_5_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_5_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_5_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_5_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42402),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23328),
            .ce(),
            .sr(N__52046));
    defparam \delay_measurement_inst.stop_timer_hc_LC_5_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_5_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_5_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42403),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23328),
            .ce(),
            .sr(N__52046));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23618),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52472),
            .ce(),
            .sr(N__51971));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_7_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_7_12_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_7_12_3  (
            .in0(N__24276),
            .in1(N__24810),
            .in2(_gnd_net_),
            .in3(N__24534),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_7_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_7_12_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_7_12_5  (
            .in0(N__24099),
            .in1(N__24840),
            .in2(_gnd_net_),
            .in3(N__24533),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_7_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_7_12_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_7_12_7  (
            .in0(N__24759),
            .in1(N__24240),
            .in2(_gnd_net_),
            .in3(N__24535),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_13_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_13_2  (
            .in0(N__34236),
            .in1(N__32106),
            .in2(N__34786),
            .in3(N__29826),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_14_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_14_4  (
            .in0(N__24536),
            .in1(N__25113),
            .in2(_gnd_net_),
            .in3(N__24297),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_7_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_7_15_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_7_15_0  (
            .in0(N__24558),
            .in1(N__24357),
            .in2(_gnd_net_),
            .in3(N__24936),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_7_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_7_15_1 .LUT_INIT=16'b0101001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_7_15_1  (
            .in0(N__24204),
            .in1(N__25011),
            .in2(N__24580),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_7_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_7_15_6 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_7_15_6  (
            .in0(N__24231),
            .in1(N__24540),
            .in2(_gnd_net_),
            .in3(N__24732),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23778),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__51996));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23748),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__51996));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_7_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23724),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__51996));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_7_17_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_7_17_0  (
            .in0(N__34787),
            .in1(N__34258),
            .in2(N__32352),
            .in3(N__29576),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_7_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_7_17_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_7_17_2  (
            .in0(N__24475),
            .in1(N__24219),
            .in2(_gnd_net_),
            .in3(N__25026),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_7_17_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_7_17_3  (
            .in0(N__24455),
            .in1(N__24705),
            .in2(_gnd_net_),
            .in3(N__24018),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_7_17_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_7_17_4  (
            .in0(N__24033),
            .in1(N__24717),
            .in2(_gnd_net_),
            .in3(N__24454),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_7_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_7_17_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_7_17_5  (
            .in0(N__24456),
            .in1(N__24177),
            .in2(_gnd_net_),
            .in3(N__24678),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_7_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_7_17_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_7_17_6  (
            .in0(N__24666),
            .in1(N__24162),
            .in2(_gnd_net_),
            .in3(N__24457),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_7_17_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_7_17_7  (
            .in0(N__24458),
            .in1(N__24396),
            .in2(_gnd_net_),
            .in3(N__24978),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__37041),
            .in2(_gnd_net_),
            .in3(N__36970),
            .lcout(\phase_controller_inst1.stoper_tr.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_18_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_18_5  (
            .in0(N__34259),
            .in1(N__29921),
            .in2(N__34851),
            .in3(N__32204),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23916),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52426),
            .ce(),
            .sr(N__52018));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_7_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23886),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52426),
            .ce(),
            .sr(N__52018));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_19_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_7_19_3  (
            .in0(N__23862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52426),
            .ce(),
            .sr(N__52018));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_7_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23838),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52426),
            .ce(),
            .sr(N__52018));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23808),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52426),
            .ce(),
            .sr(N__52018));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_7_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_7_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_7_20_3  (
            .in0(N__34242),
            .in1(N__27293),
            .in2(N__34848),
            .in3(N__29499),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_7_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_7_20_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_7_20_7  (
            .in0(N__34243),
            .in1(N__27677),
            .in2(N__34847),
            .in3(N__29742),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_7_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_7_21_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_7_21_0  (
            .in0(N__34260),
            .in1(N__34772),
            .in2(N__27227),
            .in3(N__29457),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_7_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_7_21_4 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_7_21_4  (
            .in0(N__27608),
            .in1(N__29700),
            .in2(N__34266),
            .in3(N__34773),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_7_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_7_21_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_7_21_7  (
            .in0(N__34774),
            .in1(N__34264),
            .in2(N__29580),
            .in3(N__32345),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_7_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_7_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_7_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23991),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52409),
            .ce(),
            .sr(N__52037));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_22_7 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_7_22_7  (
            .in0(N__44428),
            .in1(N__42413),
            .in2(_gnd_net_),
            .in3(N__44335),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52409),
            .ce(),
            .sr(N__52037));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_7_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_7_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_7_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52634),
            .lcout(pwm_duty_input_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52404),
            .ce(),
            .sr(N__52042));
    defparam \phase_controller_inst2.state_2_LC_8_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_8_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_8_5_0 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst2.state_2_LC_8_5_0  (
            .in0(N__28061),
            .in1(N__25841),
            .in2(N__23957),
            .in3(N__25802),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52496),
            .ce(),
            .sr(N__51941));
    defparam \phase_controller_inst2.start_timer_hc_LC_8_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_8_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_8_5_4 .LUT_INIT=16'b1100110011111000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_8_5_4  (
            .in0(N__23950),
            .in1(N__25840),
            .in2(N__32797),
            .in3(N__25801),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52496),
            .ce(),
            .sr(N__51941));
    defparam \phase_controller_inst2.state_1_LC_8_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_8_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_8_5_5 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \phase_controller_inst2.state_1_LC_8_5_5  (
            .in0(N__25272),
            .in1(N__28062),
            .in2(N__25803),
            .in3(N__25240),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52496),
            .ce(),
            .sr(N__51941));
    defparam \phase_controller_inst2.state_RNO_0_3_LC_8_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_8_6_3 .LUT_INIT=16'b0010101000111111;
    LogicCell40 \phase_controller_inst2.state_RNO_0_3_LC_8_6_3  (
            .in0(N__23961),
            .in1(N__25196),
            .in2(N__25218),
            .in3(N__25831),
            .lcout(\phase_controller_inst2.state_ns_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_flag_LC_8_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_flag_LC_8_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_flag_LC_8_7_1 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \phase_controller_inst2.start_flag_LC_8_7_1  (
            .in0(N__36565),
            .in1(N__24070),
            .in2(N__24059),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52487),
            .ce(),
            .sr(N__51947));
    defparam \phase_controller_inst2.state_4_LC_8_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_4_LC_8_7_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst2.state_4_LC_8_7_3 .LUT_INIT=16'b1100010011000100;
    LogicCell40 \phase_controller_inst2.state_4_LC_8_7_3  (
            .in0(N__36567),
            .in1(N__24072),
            .in2(N__24060),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52487),
            .ce(),
            .sr(N__51947));
    defparam \phase_controller_inst2.state_3_LC_8_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_8_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_8_7_7 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \phase_controller_inst2.state_3_LC_8_7_7  (
            .in0(N__36566),
            .in1(N__24071),
            .in2(N__24058),
            .in3(N__24039),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52487),
            .ce(),
            .sr(N__51947));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__25062),
            .in2(N__25344),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_11_1  (
            .in0(N__29879),
            .in1(N__25656),
            .in2(N__25164),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__34446),
            .in2(N__26424),
            .in3(N__29880),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__25350),
            .in2(N__34637),
            .in3(N__24021),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__34450),
            .in2(N__26358),
            .in3(N__24006),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__25176),
            .in2(N__34638),
            .in3(N__24180),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__34454),
            .in2(N__25386),
            .in3(N__24165),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__25155),
            .in2(N__34639),
            .in3(N__24150),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__34458),
            .in2(N__26316),
            .in3(N__24138),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__25329),
            .in2(N__34640),
            .in3(N__24126),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__34462),
            .in2(N__25323),
            .in3(N__24114),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__25314),
            .in2(N__34641),
            .in3(N__24102),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__34466),
            .in2(N__25308),
            .in3(N__24093),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__25170),
            .in2(N__34642),
            .in3(N__24075),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__34470),
            .in2(N__26340),
            .in3(N__24270),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__28569),
            .in2(N__34643),
            .in3(N__24255),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__34580),
            .in2(N__25443),
            .in3(N__24243),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__25335),
            .in2(N__34743),
            .in3(N__24234),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__34584),
            .in2(N__25299),
            .in3(N__24222),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__25431),
            .in2(N__34744),
            .in3(N__24207),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__34588),
            .in2(N__26520),
            .in3(N__24195),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__25290),
            .in2(N__34745),
            .in3(N__24183),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__34592),
            .in2(N__24405),
            .in3(N__24384),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__25563),
            .in2(N__34746),
            .in3(N__24372),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__34613),
            .in2(N__24369),
            .in3(N__24351),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__25404),
            .in2(N__34763),
            .in3(N__24339),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__34617),
            .in2(N__26583),
            .in3(N__24327),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__26325),
            .in2(N__34764),
            .in3(N__24312),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__34621),
            .in2(N__25425),
            .in3(N__24300),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__25503),
            .in2(N__34765),
            .in3(N__24291),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__25509),
            .in2(N__34785),
            .in3(N__24420),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_14_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_14_7  (
            .in0(N__29031),
            .in1(N__25077),
            .in2(N__24579),
            .in3(N__24417),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_8_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__29012),
            .in2(N__29881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_8_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__46342),
            .in2(N__25371),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_8_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__46346),
            .in2(N__26436),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_8_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__46343),
            .in2(N__26478),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_8_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__46347),
            .in2(N__26448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_8_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__46344),
            .in2(N__26463),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_8_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__46348),
            .in2(N__25413),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_8_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__46345),
            .in2(N__25359),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_8_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__46361),
            .in2(N__26532),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_8_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_8_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__25497),
            .in2(N__46481),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_8_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_8_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__46349),
            .in2(N__26490),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_8_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_8_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__25449),
            .in2(N__46478),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_8_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_8_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__46353),
            .in2(N__25458),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_8_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_8_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__25491),
            .in2(N__46479),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_8_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_8_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__46357),
            .in2(N__26502),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_8_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_8_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__25464),
            .in2(N__46480),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__25485),
            .in2(N__46482),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_8_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__46368),
            .in2(N__25536),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_8_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__25551),
            .in2(N__46483),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_8_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__46372),
            .in2(N__25545),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_8_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__25575),
            .in2(N__46484),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_8_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__46376),
            .in2(N__25527),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_8_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__25569),
            .in2(N__46485),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_8_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__46380),
            .in2(N__25584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_8_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__46381),
            .in2(N__26673),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_8_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__25608),
            .in2(N__46486),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_8_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__46385),
            .in2(N__26568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_8_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__26661),
            .in2(N__46487),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_8_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__46389),
            .in2(N__25680),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_8_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__25686),
            .in2(N__46488),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_8_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__46393),
            .in2(N__33711),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_8_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_8_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__34254),
            .in2(_gnd_net_),
            .in3(N__24597),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_8_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__25058),
            .in2(N__26399),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_8_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__25661),
            .in2(N__25632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_8_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__34538),
            .in2(N__25617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_8_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__25398),
            .in2(N__34733),
            .in3(N__24708),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_8_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__34542),
            .in2(N__26610),
            .in3(N__24696),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_8_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__25623),
            .in2(N__34734),
            .in3(N__24681),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__34546),
            .in2(N__25518),
            .in3(N__24669),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__26373),
            .in2(N__34735),
            .in3(N__24657),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_8_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__34550),
            .in2(N__33393),
            .in3(N__24642),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__34551),
            .in2(N__25602),
            .in3(N__24624),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__24621),
            .in2(N__34736),
            .in3(N__24600),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__34555),
            .in2(N__24867),
            .in3(N__24843),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_8_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__33612),
            .in2(N__34737),
            .in3(N__24828),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_8_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__34559),
            .in2(N__33207),
            .in3(N__24813),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_8_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_8_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__26544),
            .in2(N__34738),
            .in3(N__24795),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_8_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_8_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(N__34563),
            .in2(N__33303),
            .in3(N__24777),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_8_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(N__34564),
            .in2(N__25479),
            .in3(N__24762),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_8_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(N__26556),
            .in2(N__34739),
            .in3(N__24744),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_8_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(N__34568),
            .in2(N__24741),
            .in3(N__24720),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_8_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(N__25035),
            .in2(N__34740),
            .in3(N__25014),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_8_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_8_21_4  (
            .in0(_gnd_net_),
            .in1(N__34572),
            .in2(N__26625),
            .in3(N__24999),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_8_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_8_21_5  (
            .in0(_gnd_net_),
            .in1(N__27027),
            .in2(N__34741),
            .in3(N__24981),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_8_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_8_21_6  (
            .in0(_gnd_net_),
            .in1(N__34576),
            .in2(N__29799),
            .in3(N__24966),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_8_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(N__33861),
            .in2(N__34742),
            .in3(N__24945),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_8_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(N__24942),
            .in2(N__34843),
            .in3(N__24924),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_8_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(N__34750),
            .in2(N__26598),
            .in3(N__24906),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_8_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__33492),
            .in2(N__34844),
            .in3(N__24885),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_8_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(N__34754),
            .in2(N__26640),
            .in3(N__25149),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_8_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(N__26652),
            .in2(N__34845),
            .in3(N__25131),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_8_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_8_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(N__34758),
            .in2(N__25128),
            .in3(N__25101),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_8_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_8_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_8_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_8_22_6  (
            .in0(_gnd_net_),
            .in1(N__29838),
            .in2(N__34846),
            .in3(N__25083),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_8_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_8_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_8_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_8_22_7  (
            .in0(N__34265),
            .in1(N__34762),
            .in2(_gnd_net_),
            .in3(N__25080),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_23_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_23_4  (
            .in0(N__46489),
            .in1(N__25980),
            .in2(_gnd_net_),
            .in3(N__29019),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_23_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_23_5  (
            .in0(N__26400),
            .in1(_gnd_net_),
            .in2(N__25065),
            .in3(N__46490),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_8_26_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_26_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25284),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52387),
            .ce(),
            .sr(N__52047));
    defparam \phase_controller_inst2.start_timer_tr_LC_9_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_9_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_9_5_7 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_9_5_7  (
            .in0(N__25241),
            .in1(N__25779),
            .in2(N__25280),
            .in3(N__28033),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52493),
            .ce(),
            .sr(N__51935));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_9_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_9_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_9_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28028),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52488),
            .ce(),
            .sr(N__51942));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_9_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_9_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_9_6_4 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_9_6_4  (
            .in0(N__25216),
            .in1(N__27990),
            .in2(N__25185),
            .in3(N__28731),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52488),
            .ce(),
            .sr(N__51942));
    defparam \phase_controller_inst2.state_0_LC_9_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_9_6_7 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst2.state_0_LC_9_6_7  (
            .in0(N__25273),
            .in1(N__25248),
            .in2(N__25200),
            .in3(N__25217),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52488),
            .ce(),
            .sr(N__51942));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_9_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_9_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__28766),
            .in2(_gnd_net_),
            .in3(N__28034),
            .lcout(\phase_controller_inst2.stoper_tr.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_9_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_9_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28776),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_9_10_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_9_10_7  (
            .in0(N__28416),
            .in1(N__28396),
            .in2(_gnd_net_),
            .in3(N__28378),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_12_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_12_0  (
            .in0(N__34065),
            .in1(N__34491),
            .in2(N__26865),
            .in3(N__29159),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_9_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_9_12_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_9_12_2  (
            .in0(N__34067),
            .in1(N__34493),
            .in2(N__33255),
            .in3(N__33285),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_12_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_12_3  (
            .in0(N__33161),
            .in1(N__34063),
            .in2(N__29310),
            .in3(N__25657),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_9_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_9_12_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_9_12_4  (
            .in0(N__34066),
            .in1(N__34492),
            .in2(N__26739),
            .in3(N__29088),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_12_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_12_5  (
            .in0(N__34490),
            .in1(N__34064),
            .in2(N__29238),
            .in3(N__26976),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_9_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_9_12_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_9_12_6  (
            .in0(N__34062),
            .in1(N__26409),
            .in2(_gnd_net_),
            .in3(N__28809),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_13_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_13_1  (
            .in0(N__34077),
            .in1(N__27738),
            .in2(N__34793),
            .in3(N__29778),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_13_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_13_3  (
            .in0(N__34073),
            .in1(N__27354),
            .in2(N__34791),
            .in3(N__29535),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_13_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_13_4  (
            .in0(N__29498),
            .in1(N__34676),
            .in2(N__27294),
            .in3(N__34074),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_13_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_13_5  (
            .in0(N__34075),
            .in1(N__34681),
            .in2(N__27228),
            .in3(N__29456),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_9_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_9_13_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_9_13_6  (
            .in0(N__33642),
            .in1(N__34677),
            .in2(N__33690),
            .in3(N__34076),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_9_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_9_13_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_9_13_7  (
            .in0(N__34078),
            .in1(N__27678),
            .in2(N__34792),
            .in3(N__29738),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_14_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_14_0  (
            .in0(N__34683),
            .in1(N__34088),
            .in2(N__27489),
            .in3(N__29618),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_1  (
            .in0(N__34086),
            .in1(N__34685),
            .in2(N__32157),
            .in3(N__29361),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_9_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_9_14_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_9_14_3  (
            .in0(N__34087),
            .in1(N__34684),
            .in2(N__27612),
            .in3(N__29699),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_14_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_14_4  (
            .in0(N__34682),
            .in1(N__34089),
            .in2(N__33600),
            .in3(N__29952),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_9_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_9_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_9_15_0  (
            .in0(N__28944),
            .in1(N__26799),
            .in2(_gnd_net_),
            .in3(N__29113),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_9_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_9_15_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_9_15_1  (
            .in0(N__32301),
            .in1(N__34135),
            .in2(N__30030),
            .in3(N__34799),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_15_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_15_2  (
            .in0(N__34133),
            .in1(N__26972),
            .in2(N__34852),
            .in3(N__29231),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_9_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_9_15_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_9_15_3  (
            .in0(N__29114),
            .in1(N__34134),
            .in2(N__26805),
            .in3(N__34797),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_15_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_15_4  (
            .in0(N__28943),
            .in1(N__29299),
            .in2(_gnd_net_),
            .in3(N__33154),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_9_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_9_15_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_9_15_5  (
            .in0(N__26730),
            .in1(N__28945),
            .in2(_gnd_net_),
            .in3(N__29083),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_9_15_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_9_15_6  (
            .in0(N__34800),
            .in1(N__34235),
            .in2(N__29889),
            .in3(N__33729),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_9_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_9_15_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_9_15_7  (
            .in0(N__34234),
            .in1(N__34798),
            .in2(N__32211),
            .in3(N__29922),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_16_0  (
            .in0(N__28946),
            .in1(N__27346),
            .in2(_gnd_net_),
            .in3(N__29527),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_9_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_9_16_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_9_16_1  (
            .in0(N__33241),
            .in1(N__33280),
            .in2(_gnd_net_),
            .in3(N__28949),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_16_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_16_2  (
            .in0(N__28951),
            .in1(N__29356),
            .in2(_gnd_net_),
            .in3(N__32149),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_9_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_9_16_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_9_16_4  (
            .in0(N__34229),
            .in1(N__29357),
            .in2(N__34853),
            .in3(N__32150),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_9_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_9_16_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_9_16_5  (
            .in0(N__33328),
            .in1(N__28950),
            .in2(_gnd_net_),
            .in3(N__33367),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_16_6  (
            .in0(N__28948),
            .in1(N__33682),
            .in2(_gnd_net_),
            .in3(N__33637),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_9_16_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_9_16_7  (
            .in0(N__27226),
            .in1(N__28947),
            .in2(_gnd_net_),
            .in3(N__29446),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_17_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_17_0  (
            .in0(N__33916),
            .in1(N__28958),
            .in2(_gnd_net_),
            .in3(N__33880),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_9_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_9_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_9_17_1  (
            .in0(N__28956),
            .in1(N__27546),
            .in2(_gnd_net_),
            .in3(N__29650),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_9_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_9_17_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_9_17_2  (
            .in0(N__29822),
            .in1(N__28957),
            .in2(_gnd_net_),
            .in3(N__32102),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_3  (
            .in0(N__33881),
            .in1(N__34230),
            .in2(N__34854),
            .in3(N__33917),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_17_4  (
            .in0(N__28953),
            .in1(N__27673),
            .in2(_gnd_net_),
            .in3(N__29731),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_9_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_9_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_9_17_5  (
            .in0(N__28955),
            .in1(N__27604),
            .in2(_gnd_net_),
            .in3(N__29689),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_9_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_9_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_9_17_6  (
            .in0(N__28952),
            .in1(N__27734),
            .in2(_gnd_net_),
            .in3(N__29774),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_17_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_17_7  (
            .in0(N__27482),
            .in1(N__29611),
            .in2(_gnd_net_),
            .in3(N__28954),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_18_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_18_0  (
            .in0(N__34809),
            .in1(N__34195),
            .in2(N__26803),
            .in3(N__29118),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_18_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_18_1  (
            .in0(N__34191),
            .in1(N__29917),
            .in2(_gnd_net_),
            .in3(N__32197),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_18_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_18_2  (
            .in0(N__33589),
            .in1(N__34190),
            .in2(_gnd_net_),
            .in3(N__29945),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_18_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_18_3  (
            .in0(N__34192),
            .in1(N__29309),
            .in2(N__25671),
            .in3(N__33162),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_18_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_18_4  (
            .in0(N__34808),
            .in1(N__34194),
            .in2(N__29160),
            .in3(N__26861),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_9_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_9_18_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_9_18_5  (
            .in0(N__34193),
            .in1(N__34810),
            .in2(N__27015),
            .in3(N__29274),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_18_6  (
            .in0(N__32293),
            .in1(N__34189),
            .in2(_gnd_net_),
            .in3(N__30023),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_18_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_18_7  (
            .in0(N__34196),
            .in1(N__34807),
            .in2(N__27353),
            .in3(N__29534),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_9_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_9_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_9_19_0  (
            .in0(N__25969),
            .in1(N__28828),
            .in2(_gnd_net_),
            .in3(N__25590),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_1_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_9_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_9_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_9_19_1  (
            .in0(N__25957),
            .in1(N__33181),
            .in2(_gnd_net_),
            .in3(N__25587),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_2_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_9_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_9_19_2  (
            .in0(N__25970),
            .in1(N__26939),
            .in2(_gnd_net_),
            .in3(N__25713),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_3_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_9_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_9_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_9_19_3  (
            .in0(N__25958),
            .in1(N__26885),
            .in2(_gnd_net_),
            .in3(N__25710),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_4_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_9_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_9_19_4  (
            .in0(N__25971),
            .in1(N__26825),
            .in2(_gnd_net_),
            .in3(N__25707),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_5_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_9_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_9_19_5  (
            .in0(N__25959),
            .in1(N__26759),
            .in2(_gnd_net_),
            .in3(N__25704),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_6_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_9_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_9_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_9_19_6  (
            .in0(N__25972),
            .in1(N__26696),
            .in2(_gnd_net_),
            .in3(N__25701),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_7_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_9_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_9_19_7  (
            .in0(N__25960),
            .in1(N__27374),
            .in2(_gnd_net_),
            .in3(N__25698),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__52415),
            .ce(N__32610),
            .sr(N__52002));
    defparam \current_shift_inst.timer_s1.counter_8_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_9_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_9_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_9_20_0  (
            .in0(N__25956),
            .in1(N__27314),
            .in2(_gnd_net_),
            .in3(N__25695),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_9_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_9_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_9_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_9_20_1  (
            .in0(N__25968),
            .in1(N__27248),
            .in2(_gnd_net_),
            .in3(N__25692),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_10_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_9_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_9_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_9_20_2  (
            .in0(N__25953),
            .in1(N__27179),
            .in2(_gnd_net_),
            .in3(N__25689),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_11_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_9_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_9_20_3  (
            .in0(N__25965),
            .in1(N__27155),
            .in2(_gnd_net_),
            .in3(N__25740),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_12_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_9_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_9_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_9_20_4  (
            .in0(N__25954),
            .in1(N__27131),
            .in2(_gnd_net_),
            .in3(N__25737),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_13_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_9_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_9_20_5  (
            .in0(N__25966),
            .in1(N__27074),
            .in2(_gnd_net_),
            .in3(N__25734),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_14_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_9_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_9_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_9_20_6  (
            .in0(N__25955),
            .in1(N__27050),
            .in2(_gnd_net_),
            .in3(N__25731),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_15_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_9_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_9_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_9_20_7  (
            .in0(N__25967),
            .in1(N__27758),
            .in2(_gnd_net_),
            .in3(N__25728),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__52410),
            .ce(N__32609),
            .sr(N__52010));
    defparam \current_shift_inst.timer_s1.counter_16_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_9_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_9_21_0  (
            .in0(N__25944),
            .in1(N__27698),
            .in2(_gnd_net_),
            .in3(N__25725),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_17_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_9_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_9_21_1  (
            .in0(N__25961),
            .in1(N__27632),
            .in2(_gnd_net_),
            .in3(N__25722),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_18_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_9_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_9_21_2  (
            .in0(N__25945),
            .in1(N__27566),
            .in2(_gnd_net_),
            .in3(N__25719),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_19_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_9_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_9_21_3  (
            .in0(N__25962),
            .in1(N__27509),
            .in2(_gnd_net_),
            .in3(N__25716),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_20_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_9_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_9_21_4  (
            .in0(N__25946),
            .in1(N__27446),
            .in2(_gnd_net_),
            .in3(N__25770),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_21_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_9_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_9_21_5  (
            .in0(N__25963),
            .in1(N__27422),
            .in2(_gnd_net_),
            .in3(N__25767),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_22_LC_9_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_9_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_9_21_6  (
            .in0(N__25947),
            .in1(N__27398),
            .in2(_gnd_net_),
            .in3(N__25764),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_23_LC_9_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_9_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_9_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_9_21_7  (
            .in0(N__25964),
            .in1(N__27905),
            .in2(_gnd_net_),
            .in3(N__25761),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__52405),
            .ce(N__32598),
            .sr(N__52019));
    defparam \current_shift_inst.timer_s1.counter_24_LC_9_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_9_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_9_22_0  (
            .in0(N__25931),
            .in1(N__27881),
            .in2(_gnd_net_),
            .in3(N__25758),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__52400),
            .ce(N__32602),
            .sr(N__52026));
    defparam \current_shift_inst.timer_s1.counter_25_LC_9_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_9_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_9_22_1  (
            .in0(N__25973),
            .in1(N__27857),
            .in2(_gnd_net_),
            .in3(N__25755),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__52400),
            .ce(N__32602),
            .sr(N__52026));
    defparam \current_shift_inst.timer_s1.counter_26_LC_9_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_9_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_9_22_2  (
            .in0(N__25932),
            .in1(N__27821),
            .in2(_gnd_net_),
            .in3(N__25752),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__52400),
            .ce(N__32602),
            .sr(N__52026));
    defparam \current_shift_inst.timer_s1.counter_27_LC_9_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_9_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_9_22_3  (
            .in0(N__25974),
            .in1(N__27785),
            .in2(_gnd_net_),
            .in3(N__25749),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__52400),
            .ce(N__32602),
            .sr(N__52026));
    defparam \current_shift_inst.timer_s1.counter_28_LC_9_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_9_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_9_22_4  (
            .in0(N__25933),
            .in1(N__27834),
            .in2(_gnd_net_),
            .in3(N__25746),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__52400),
            .ce(N__32602),
            .sr(N__52026));
    defparam \current_shift_inst.timer_s1.counter_29_LC_9_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_9_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_9_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_9_22_5  (
            .in0(N__27798),
            .in1(N__25934),
            .in2(_gnd_net_),
            .in3(N__25743),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52400),
            .ce(N__32602),
            .sr(N__52026));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_9_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_9_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_9_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28981),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52396),
            .ce(N__33754),
            .sr(N__52033));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_9_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_9_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33529),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40929),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_27_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25845),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52379),
            .ce(),
            .sr(N__52048));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_5_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_5_0  (
            .in0(N__25797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28051),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_10_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_10_6_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_10_6_5  (
            .in0(N__28027),
            .in1(N__52083),
            .in2(_gnd_net_),
            .in3(N__28765),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__32802),
            .in2(_gnd_net_),
            .in3(N__38215),
            .lcout(\phase_controller_inst2.stoper_hc.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_10_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_10_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_0_LC_10_7_0  (
            .in0(N__26284),
            .in1(N__27969),
            .in2(N__28703),
            .in3(N__28704),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_0 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_10_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_10_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_1_LC_10_7_1  (
            .in0(N__26292),
            .in1(N__27948),
            .in2(_gnd_net_),
            .in3(N__25773),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_1 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_10_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_10_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_10_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_2_LC_10_7_2  (
            .in0(N__26285),
            .in1(N__27927),
            .in2(_gnd_net_),
            .in3(N__26007),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_2 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_10_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_10_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_3_LC_10_7_3  (
            .in0(N__26293),
            .in1(N__28251),
            .in2(_gnd_net_),
            .in3(N__26004),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_3 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_10_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_10_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_4_LC_10_7_4  (
            .in0(N__26286),
            .in1(N__28230),
            .in2(_gnd_net_),
            .in3(N__26001),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_4 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_10_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_10_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_5_LC_10_7_5  (
            .in0(N__26294),
            .in1(N__28209),
            .in2(_gnd_net_),
            .in3(N__25998),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_5 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_10_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_10_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_6_LC_10_7_6  (
            .in0(N__26287),
            .in1(N__28188),
            .in2(_gnd_net_),
            .in3(N__25995),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_6 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_10_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_10_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_10_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_7_LC_10_7_7  (
            .in0(N__26295),
            .in1(N__28167),
            .in2(_gnd_net_),
            .in3(N__25992),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_7 ),
            .clk(N__52473),
            .ce(N__26166),
            .sr(N__51939));
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_10_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_10_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_8_LC_10_8_0  (
            .in0(N__26283),
            .in1(N__28146),
            .in2(_gnd_net_),
            .in3(N__25989),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_8 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_10_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_10_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_10_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_9_LC_10_8_1  (
            .in0(N__26291),
            .in1(N__28125),
            .in2(_gnd_net_),
            .in3(N__25986),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_9 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_10_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_10_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_10_LC_10_8_2  (
            .in0(N__26280),
            .in1(N__28104),
            .in2(_gnd_net_),
            .in3(N__25983),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_10 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_10_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_10_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_11_LC_10_8_3  (
            .in0(N__26288),
            .in1(N__28356),
            .in2(_gnd_net_),
            .in3(N__26034),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_11 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_10_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_10_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_12_LC_10_8_4  (
            .in0(N__26281),
            .in1(N__28335),
            .in2(_gnd_net_),
            .in3(N__26031),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_12 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_10_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_10_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_10_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_13_LC_10_8_5  (
            .in0(N__26289),
            .in1(N__28314),
            .in2(_gnd_net_),
            .in3(N__26028),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_13 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_10_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_10_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_14_LC_10_8_6  (
            .in0(N__26282),
            .in1(N__28293),
            .in2(_gnd_net_),
            .in3(N__26025),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_14 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_10_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_10_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_10_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_15_LC_10_8_7  (
            .in0(N__26290),
            .in1(N__28272),
            .in2(_gnd_net_),
            .in3(N__26022),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_15 ),
            .clk(N__52466),
            .ce(N__26167),
            .sr(N__51943));
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_10_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_10_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_16_LC_10_9_0  (
            .in0(N__26272),
            .in1(N__28630),
            .in2(_gnd_net_),
            .in3(N__26019),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_16 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_10_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_10_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_17_LC_10_9_1  (
            .in0(N__26276),
            .in1(N__28606),
            .in2(_gnd_net_),
            .in3(N__26016),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_17 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_10_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_10_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_18_LC_10_9_2  (
            .in0(N__26273),
            .in1(N__28558),
            .in2(_gnd_net_),
            .in3(N__26013),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_18 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_10_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_10_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_19_LC_10_9_3  (
            .in0(N__26277),
            .in1(N__28540),
            .in2(_gnd_net_),
            .in3(N__26010),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_19 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_10_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_10_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_20_LC_10_9_4  (
            .in0(N__26274),
            .in1(N__32695),
            .in2(_gnd_net_),
            .in3(N__26061),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_20 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_10_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_10_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_21_LC_10_9_5  (
            .in0(N__26278),
            .in1(N__32713),
            .in2(_gnd_net_),
            .in3(N__26058),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_21 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_10_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_10_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_22_LC_10_9_6  (
            .in0(N__26275),
            .in1(N__32955),
            .in2(_gnd_net_),
            .in3(N__26055),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_22 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_10_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_10_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_23_LC_10_9_7  (
            .in0(N__26279),
            .in1(N__32973),
            .in2(_gnd_net_),
            .in3(N__26052),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_23 ),
            .clk(N__52461),
            .ce(N__26168),
            .sr(N__51945));
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_10_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_10_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_24_LC_10_10_0  (
            .in0(N__26264),
            .in1(N__28665),
            .in2(_gnd_net_),
            .in3(N__26049),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_24 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_10_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_10_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_25_LC_10_10_1  (
            .in0(N__26268),
            .in1(N__28680),
            .in2(_gnd_net_),
            .in3(N__26046),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_25 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_10_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_10_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_26_LC_10_10_2  (
            .in0(N__26265),
            .in1(N__32842),
            .in2(_gnd_net_),
            .in3(N__26043),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_26 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_10_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_10_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_27_LC_10_10_3  (
            .in0(N__26269),
            .in1(N__32872),
            .in2(_gnd_net_),
            .in3(N__26040),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_27 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_10_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_10_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_28_LC_10_10_4  (
            .in0(N__26266),
            .in1(N__28380),
            .in2(_gnd_net_),
            .in3(N__26037),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_28 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_10_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_10_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_29_LC_10_10_5  (
            .in0(N__26270),
            .in1(N__28398),
            .in2(_gnd_net_),
            .in3(N__26301),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_29 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_10_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_10_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_30_LC_10_10_6  (
            .in0(N__26267),
            .in1(N__28452),
            .in2(_gnd_net_),
            .in3(N__26298),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_29 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_30 ),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_10_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_31_LC_10_10_7  (
            .in0(N__26271),
            .in1(N__28470),
            .in2(_gnd_net_),
            .in3(N__26172),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52457),
            .ce(N__26169),
            .sr(N__51951));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_28_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40470),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52451),
            .ce(N__36325),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_10_11_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_10_11_2  (
            .in0(N__28468),
            .in1(N__28450),
            .in2(_gnd_net_),
            .in3(N__28419),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_10_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_10_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26151),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52444),
            .ce(),
            .sr(N__51956));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_10_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26121),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52444),
            .ce(),
            .sr(N__51956));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_10_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_10_12_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__26102),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52444),
            .ce(),
            .sr(N__51956));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_10_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_10_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26081),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52444),
            .ce(),
            .sr(N__51956));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_13_2  (
            .in0(N__28988),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52438),
            .ce(N__33759),
            .sr(N__51960));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_10_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_10_13_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_10_13_3  (
            .in0(N__27007),
            .in1(N__34061),
            .in2(N__34860),
            .in3(N__29270),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_10_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_10_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29330),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_10_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_10_13_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__34060),
            .in2(N__26403),
            .in3(N__28802),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_14_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_14_1  (
            .in0(N__26735),
            .in1(N__34068),
            .in2(N__29087),
            .in3(N__34782),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_14_2  (
            .in0(N__34069),
            .in1(N__26918),
            .in2(N__34850),
            .in3(N__29189),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_10_14_3 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_10_14_3  (
            .in0(N__29394),
            .in1(N__34784),
            .in2(N__27111),
            .in3(N__34071),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_14_4  (
            .in0(N__34072),
            .in1(N__32256),
            .in2(N__34849),
            .in3(N__29982),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_14_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_14_5  (
            .in0(N__33411),
            .in1(N__34783),
            .in2(N__33452),
            .in3(N__34070),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26856),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26734),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_0  (
            .in0(N__28881),
            .in1(N__26965),
            .in2(_gnd_net_),
            .in3(N__29224),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_1  (
            .in0(N__28883),
            .in1(N__26857),
            .in2(_gnd_net_),
            .in3(N__29143),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26964),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_3  (
            .in0(N__28882),
            .in1(N__26917),
            .in2(_gnd_net_),
            .in3(N__29185),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26804),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_10_15_5  (
            .in0(N__27279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_6  (
            .in0(N__28880),
            .in1(N__27014),
            .in2(_gnd_net_),
            .in3(N__29263),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_10_15_7  (
            .in0(N__33438),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_16_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_16_0  (
            .in0(N__34136),
            .in1(N__34893),
            .in2(N__27110),
            .in3(N__29390),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_16_1  (
            .in0(N__28908),
            .in1(N__33439),
            .in2(_gnd_net_),
            .in3(N__33409),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26916),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_10_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_10_16_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_10_16_3  (
            .in0(N__29658),
            .in1(N__34137),
            .in2(N__34908),
            .in3(N__27541),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4  (
            .in0(N__27103),
            .in1(N__28910),
            .in2(_gnd_net_),
            .in3(N__29389),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_5  (
            .in0(N__28909),
            .in1(_gnd_net_),
            .in2(N__27289),
            .in3(N__29482),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27006),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_10_16_7  (
            .in0(N__33231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_10_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_10_17_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__47157),
            .in2(_gnd_net_),
            .in3(N__47642),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52416),
            .ce(N__43466),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27603),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_10_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27213),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27540),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33669),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27474),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0  (
            .in0(N__34188),
            .in1(N__34898),
            .in2(N__33513),
            .in3(N__33545),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_10_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_10_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27723),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_10_18_2  (
            .in0(N__34185),
            .in1(N__33544),
            .in2(_gnd_net_),
            .in3(N__33508),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33357),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_18_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_18_4  (
            .in0(N__34187),
            .in1(N__34897),
            .in2(N__27733),
            .in3(N__29770),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27672),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_6  (
            .in0(N__28962),
            .in1(N__32338),
            .in2(_gnd_net_),
            .in3(N__29566),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_7  (
            .in0(N__32251),
            .in1(N__34186),
            .in2(_gnd_net_),
            .in3(N__29971),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_19_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_19_0  (
            .in0(N__34901),
            .in1(N__34202),
            .in2(N__33596),
            .in3(N__29944),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_10_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_10_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27094),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_19_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_19_2  (
            .in0(N__34899),
            .in1(N__34201),
            .in2(N__29978),
            .in3(N__32252),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27329),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_4  (
            .in0(N__34903),
            .in1(N__34198),
            .in2(N__29657),
            .in3(N__27545),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_19_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_19_5  (
            .in0(N__34197),
            .in1(N__34900),
            .in2(N__29199),
            .in3(N__26919),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_19_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_19_6  (
            .in0(N__34904),
            .in1(N__34200),
            .in2(N__32300),
            .in3(N__30022),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_7  (
            .in0(N__34199),
            .in1(N__34902),
            .in2(N__29619),
            .in3(N__27481),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_10_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_10_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__26935),
            .in2(N__28832),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_10_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_10_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__26881),
            .in2(N__33185),
            .in3(N__26943),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_10_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_10_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__26821),
            .in2(N__26940),
            .in3(N__26889),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_10_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_10_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_10_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__26755),
            .in2(N__26886),
            .in3(N__26829),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_10_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_10_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_10_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__26692),
            .in2(N__26826),
            .in3(N__26763),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_10_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_10_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_10_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__27370),
            .in2(N__26760),
            .in3(N__26700),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_10_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_10_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_10_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__27310),
            .in2(N__26697),
            .in3(N__26676),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_10_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_10_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_10_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__27244),
            .in2(N__27375),
            .in3(N__27318),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__52401),
            .ce(N__33756),
            .sr(N__51997));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_10_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_10_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__27175),
            .in2(N__27315),
            .in3(N__27252),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_10_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__27151),
            .in2(N__27249),
            .in3(N__27183),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_10_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__27127),
            .in2(N__27180),
            .in3(N__27159),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_10_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__27070),
            .in2(N__27156),
            .in3(N__27135),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_10_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_10_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__27046),
            .in2(N__27132),
            .in3(N__27078),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_10_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__27754),
            .in2(N__27075),
            .in3(N__27054),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_10_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_10_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__27694),
            .in2(N__27051),
            .in3(N__27030),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_10_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_10_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__27628),
            .in2(N__27759),
            .in3(N__27702),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__52397),
            .ce(N__33755),
            .sr(N__52003));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_10_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_10_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_10_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__27562),
            .in2(N__27699),
            .in3(N__27636),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_10_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_10_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_10_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__27505),
            .in2(N__27633),
            .in3(N__27570),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_10_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_10_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__27442),
            .in2(N__27567),
            .in3(N__27513),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_10_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_10_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_10_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__27418),
            .in2(N__27510),
            .in3(N__27450),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_10_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_10_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_10_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__27394),
            .in2(N__27447),
            .in3(N__27426),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_10_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_10_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__27901),
            .in2(N__27423),
            .in3(N__27402),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_10_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_10_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_10_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__27877),
            .in2(N__27399),
            .in3(N__27378),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_10_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_10_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_10_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__27853),
            .in2(N__27906),
            .in3(N__27885),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__52392),
            .ce(N__33753),
            .sr(N__52011));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_10_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_10_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_10_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__27817),
            .in2(N__27882),
            .in3(N__27861),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__52389),
            .ce(N__33752),
            .sr(N__52020));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_10_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_10_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_10_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__27781),
            .in2(N__27858),
            .in3(N__27837),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__52389),
            .ce(N__33752),
            .sr(N__52020));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_10_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_10_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__27833),
            .in2(N__27822),
            .in3(N__27801),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__52389),
            .ce(N__33752),
            .sr(N__52020));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_10_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_10_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_10_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(N__27797),
            .in2(N__27786),
            .in3(N__27765),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__52389),
            .ce(N__33752),
            .sr(N__52020));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_10_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_10_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27762),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_10_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_10_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_10_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37040),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52384),
            .ce(),
            .sr(N__52030));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_27_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36959),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_10_28_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_10_28_2 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_10_28_2  (
            .in0(N__35787),
            .in1(N__34950),
            .in2(_gnd_net_),
            .in3(N__35813),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_11_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_11_5_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_11_5_7  (
            .in0(N__27985),
            .in1(N__28029),
            .in2(_gnd_net_),
            .in3(N__28778),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_6_0 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_11_6_0  (
            .in0(N__38772),
            .in1(N__32817),
            .in2(N__28071),
            .in3(N__28055),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52474),
            .ce(),
            .sr(N__51932));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_11_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_11_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_11_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32801),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52474),
            .ce(),
            .sr(N__51932));
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_6_5 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_11_6_5  (
            .in0(N__32816),
            .in1(N__32800),
            .in2(N__38220),
            .in3(N__38771),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52474),
            .ce(),
            .sr(N__51932));
    defparam \phase_controller_inst2.stoper_tr.running_LC_11_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_11_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_11_6_7 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_11_6_7  (
            .in0(N__27989),
            .in1(N__28035),
            .in2(N__28782),
            .in3(N__28730),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52474),
            .ce(),
            .sr(N__51932));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_11_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_11_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__33054),
            .in2(N__27957),
            .in3(N__27968),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_11_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_11_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__32736),
            .in2(N__27936),
            .in3(N__27947),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_11_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_11_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__32742),
            .in2(N__27915),
            .in3(N__27926),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_11_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_11_7_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_11_7_3  (
            .in0(N__28250),
            .in1(N__32754),
            .in2(N__28239),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_11_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_11_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__32928),
            .in2(N__28218),
            .in3(N__28229),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_11_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_11_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__32748),
            .in2(N__28197),
            .in3(N__28208),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_11_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_11_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_11_7_6  (
            .in0(N__28187),
            .in1(N__33009),
            .in2(N__28176),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_11_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_11_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__36426),
            .in2(N__28155),
            .in3(N__28166),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__32730),
            .in2(N__28134),
            .in3(N__28145),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_8 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__32916),
            .in2(N__28113),
            .in3(N__28124),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_11_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_11_8_2  (
            .in0(N__28103),
            .in1(N__33066),
            .in2(N__28092),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_11_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__33042),
            .in2(N__28344),
            .in3(N__28355),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_11_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__32991),
            .in2(N__28323),
            .in3(N__28334),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_11_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_11_8_5  (
            .in0(N__28313),
            .in1(N__32907),
            .in2(N__28302),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_11_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_11_8_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_11_8_6  (
            .in0(N__28292),
            .in1(N__33480),
            .in2(N__28281),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_11_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_11_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__36489),
            .in2(N__28260),
            .in3(N__28271),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__28590),
            .in2(N__28644),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_11_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__28581),
            .in2(N__28524),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_11_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__32679),
            .in2(N__32724),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_11_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__32979),
            .in2(N__32937),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_11_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__28650),
            .in2(N__28428),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_11_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__28509),
            .in2(N__33120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_11_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__28362),
            .in2(N__28500),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_11_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__28434),
            .in2(N__28485),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28473),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_10_2 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_10_2  (
            .in0(N__28418),
            .in1(N__28469),
            .in2(_gnd_net_),
            .in3(N__28451),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_11_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_11_10_3 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_11_10_3  (
            .in0(N__28678),
            .in1(N__28663),
            .in2(N__33029),
            .in3(N__32888),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_10_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_10_4  (
            .in0(N__28417),
            .in1(N__28397),
            .in2(_gnd_net_),
            .in3(N__28379),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_11_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_11_10_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__28777),
            .in2(_gnd_net_),
            .in3(N__28720),
            .lcout(\phase_controller_inst2.stoper_tr.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_11_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_11_10_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_11_10_6  (
            .in0(N__52084),
            .in1(N__33105),
            .in2(_gnd_net_),
            .in3(N__39209),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_10_7 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_10_7  (
            .in0(N__28679),
            .in1(N__28664),
            .in2(N__33030),
            .in3(N__32889),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_11_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_11_11_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_11_11_0  (
            .in0(N__36393),
            .in1(N__28632),
            .in2(N__28614),
            .in3(N__32898),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_11_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_11_11_2 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_11_11_2  (
            .in0(N__36392),
            .in1(N__28631),
            .in2(N__28613),
            .in3(N__32897),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_11_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_11_12_0 .LUT_INIT=16'b1101010011011101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_11_12_0  (
            .in0(N__28541),
            .in1(N__36377),
            .in2(N__36411),
            .in3(N__28559),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_12_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_12_1  (
            .in0(N__34079),
            .in1(N__33378),
            .in2(N__34859),
            .in3(N__33333),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_11_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_11_12_3 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_11_12_3  (
            .in0(N__28560),
            .in1(N__36407),
            .in2(N__36378),
            .in3(N__28542),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_11_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_11_12_5 .LUT_INIT=16'b1000101011101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_11_12_5  (
            .in0(N__36477),
            .in1(N__36030),
            .in2(N__32849),
            .in3(N__32876),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__33096),
            .in2(_gnd_net_),
            .in3(N__39197),
            .lcout(\phase_controller_inst1.stoper_hc.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_11_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_11_13_2 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_11_13_2  (
            .in0(N__29043),
            .in1(N__29049),
            .in2(N__39231),
            .in3(N__36783),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52433),
            .ce(),
            .sr(N__51957));
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_13_5 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_11_13_5  (
            .in0(N__33095),
            .in1(N__29042),
            .in2(N__39207),
            .in3(N__39230),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52433),
            .ce(),
            .sr(N__51957));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_13_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_13_6  (
            .in0(N__29041),
            .in1(N__33094),
            .in2(_gnd_net_),
            .in3(N__39193),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_11_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_11_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__34090),
            .in2(_gnd_net_),
            .in3(N__34775),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28800),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_14_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_14_5  (
            .in0(N__28801),
            .in1(_gnd_net_),
            .in2(N__29022),
            .in3(N__28876),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28995),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52428),
            .ce(N__33758),
            .sr(N__51961));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28839),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52428),
            .ce(N__33758),
            .sr(N__51961));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__33459),
            .in2(N__29334),
            .in3(N__29329),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__29280),
            .in2(_gnd_net_),
            .in3(N__29247),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__29244),
            .in2(_gnd_net_),
            .in3(N__29208),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__29205),
            .in2(_gnd_net_),
            .in3(N__29169),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__29166),
            .in2(_gnd_net_),
            .in3(N__29127),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__29124),
            .in2(_gnd_net_),
            .in3(N__29097),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__29094),
            .in2(_gnd_net_),
            .in3(N__29061),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__29058),
            .in2(_gnd_net_),
            .in3(N__29052),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_16_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29547),
            .in3(N__29508),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__29505),
            .in2(_gnd_net_),
            .in3(N__29466),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__29463),
            .in2(_gnd_net_),
            .in3(N__29424),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__29421),
            .in2(_gnd_net_),
            .in3(N__29415),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__29412),
            .in2(_gnd_net_),
            .in3(N__29406),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__29403),
            .in2(_gnd_net_),
            .in3(N__29376),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__29373),
            .in2(_gnd_net_),
            .in3(N__29364),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__32121),
            .in2(_gnd_net_),
            .in3(N__29337),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__29784),
            .in2(_gnd_net_),
            .in3(N__29751),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__29748),
            .in2(_gnd_net_),
            .in3(N__29709),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__29706),
            .in2(_gnd_net_),
            .in3(N__29667),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__29664),
            .in2(_gnd_net_),
            .in3(N__29628),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__29625),
            .in2(_gnd_net_),
            .in3(N__29589),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__32064),
            .in2(_gnd_net_),
            .in3(N__29586),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__33696),
            .in2(_gnd_net_),
            .in3(N__29583),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__32310),
            .in2(_gnd_net_),
            .in3(N__29550),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__32265),
            .in2(_gnd_net_),
            .in3(N__30003),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__30000),
            .in2(_gnd_net_),
            .in3(N__29985),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__32223),
            .in2(_gnd_net_),
            .in3(N__29955),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__33555),
            .in2(_gnd_net_),
            .in3(N__29925),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__32166),
            .in2(_gnd_net_),
            .in3(N__29895),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29892),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_18_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_18_6  (
            .in0(N__29888),
            .in1(N__34887),
            .in2(N__29841),
            .in3(N__34238),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_18_7  (
            .in0(N__34237),
            .in1(N__32098),
            .in2(N__34905),
            .in3(N__29818),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_11_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_11_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__36729),
            .in2(N__36708),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_11_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_11_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__30435),
            .in2(N__30408),
            .in3(N__30393),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_11_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_11_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__30390),
            .in2(N__30375),
            .in3(N__30324),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_11_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_11_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_11_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__30321),
            .in2(N__30309),
            .in3(N__30270),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_11_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_11_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__30267),
            .in2(N__30252),
            .in3(N__30204),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_11_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_11_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_11_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__30201),
            .in2(N__30186),
            .in3(N__30147),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_11_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_11_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_11_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__30144),
            .in2(N__30129),
            .in3(N__30084),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_11_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_11_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_11_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__30081),
            .in2(N__30072),
            .in3(N__30033),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__52402),
            .ce(),
            .sr(N__51986));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_11_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_11_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_11_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__30954),
            .in2(N__30942),
            .in3(N__30894),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_11_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_11_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_11_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__30891),
            .in2(N__30873),
            .in3(N__30825),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_11_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_11_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_11_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__30822),
            .in2(N__30807),
            .in3(N__30756),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_11_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_11_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_11_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__30753),
            .in2(N__30738),
            .in3(N__30687),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_11_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_11_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_11_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__30684),
            .in2(N__30669),
            .in3(N__30627),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_11_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_11_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_11_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__30624),
            .in2(N__30609),
            .in3(N__30573),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_11_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_11_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_11_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__30570),
            .in2(N__30555),
            .in3(N__30498),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_11_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_11_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_11_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(N__30495),
            .in2(N__30483),
            .in3(N__30438),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__52398),
            .ce(),
            .sr(N__51993));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_11_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_11_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_11_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__31452),
            .in2(N__31443),
            .in3(N__31392),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_11_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_11_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_11_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__31389),
            .in2(N__31374),
            .in3(N__31329),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_11_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_11_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_11_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__31326),
            .in2(N__31308),
            .in3(N__31260),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_11_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_11_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__31257),
            .in2(N__31242),
            .in3(N__31188),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_11_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_11_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_11_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__31185),
            .in2(N__31173),
            .in3(N__31134),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_11_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_11_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_11_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__31131),
            .in2(N__31119),
            .in3(N__31077),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_11_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_11_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_11_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__31074),
            .in2(N__31062),
            .in3(N__31017),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_11_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_11_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_11_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__31014),
            .in2(N__30999),
            .in3(N__30957),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__52393),
            .ce(),
            .sr(N__51998));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_11_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_11_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_11_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__32046),
            .in2(N__32028),
            .in3(N__31983),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_11_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_11_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_11_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__31980),
            .in2(N__31965),
            .in3(N__31920),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_11_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_11_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__31917),
            .in2(N__31899),
            .in3(N__31851),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_11_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_11_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__31848),
            .in2(N__31839),
            .in3(N__31785),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_11_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_11_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_11_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__31782),
            .in2(N__31764),
            .in3(N__31725),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_11_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_11_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_11_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__31722),
            .in2(N__31713),
            .in3(N__31662),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_11_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_11_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_11_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_11_22_6  (
            .in0(N__31659),
            .in1(N__31488),
            .in2(_gnd_net_),
            .in3(N__31473),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52390),
            .ce(),
            .sr(N__52004));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_23_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_23_0  (
            .in0(N__36885),
            .in1(N__37036),
            .in2(_gnd_net_),
            .in3(N__36949),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32328),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32276),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_23_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__32234),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32182),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32140),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_11_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_11_24_1 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_11_24_1  (
            .in0(N__35844),
            .in1(N__35300),
            .in2(N__35876),
            .in3(N__35286),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_24_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__32088),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_11_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_11_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__32052),
            .in2(N__34986),
            .in3(N__35247),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_0 ),
            .ltout(),
            .carryin(bfn_11_25_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_11_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_11_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_11_25_1  (
            .in0(_gnd_net_),
            .in1(N__35082),
            .in2(N__32439),
            .in3(N__35232),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_11_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_11_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_11_25_2  (
            .in0(_gnd_net_),
            .in1(N__35076),
            .in2(N__32430),
            .in3(N__35214),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_11_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_11_25_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_11_25_3  (
            .in0(_gnd_net_),
            .in1(N__35088),
            .in2(N__32421),
            .in3(N__35193),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_11_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_11_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_11_25_4  (
            .in0(_gnd_net_),
            .in1(N__35307),
            .in2(N__32412),
            .in3(N__35172),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_11_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_11_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(N__35094),
            .in2(N__32400),
            .in3(N__35154),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_11_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_11_25_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_11_25_6  (
            .in0(N__35469),
            .in1(N__35070),
            .in2(N__32391),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_11_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_11_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(N__33813),
            .in2(N__32379),
            .in3(N__35451),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_11_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_11_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_11_26_0  (
            .in0(_gnd_net_),
            .in1(N__35064),
            .in2(N__32370),
            .in3(N__35433),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_8 ),
            .ltout(),
            .carryin(bfn_11_26_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_11_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_11_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_11_26_1  (
            .in0(_gnd_net_),
            .in1(N__35019),
            .in2(N__32361),
            .in3(N__35415),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_11_26_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_11_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_11_26_2  (
            .in0(_gnd_net_),
            .in1(N__33837),
            .in2(N__32505),
            .in3(N__35397),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_11_26_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_11_26_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__33801),
            .in2(N__32496),
            .in3(N__35379),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_11_26_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_11_26_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_11_26_4  (
            .in0(_gnd_net_),
            .in1(N__33825),
            .in2(N__32484),
            .in3(N__35361),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_11_26_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_11_26_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_11_26_5  (
            .in0(N__35343),
            .in1(N__35058),
            .in2(N__32472),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_11_26_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_11_26_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_11_26_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_11_26_6  (
            .in0(N__35325),
            .in1(N__33789),
            .in2(N__32460),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_11_26_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_11_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(N__33849),
            .in2(N__32448),
            .in3(N__35562),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_11_27_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_11_27_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_11_27_0  (
            .in0(_gnd_net_),
            .in1(N__37932),
            .in2(N__37851),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_27_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_11_27_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_11_27_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_11_27_1  (
            .in0(_gnd_net_),
            .in1(N__38283),
            .in2(N__38358),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_11_27_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_11_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_11_27_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_11_27_2  (
            .in0(_gnd_net_),
            .in1(N__32664),
            .in2(N__32652),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_11_27_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_11_27_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_11_27_3  (
            .in0(_gnd_net_),
            .in1(N__32658),
            .in2(N__32673),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_11_27_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_11_27_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_11_27_4  (
            .in0(_gnd_net_),
            .in1(N__32619),
            .in2(N__32640),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_11_27_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_11_27_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_11_27_5  (
            .in0(_gnd_net_),
            .in1(N__35268),
            .in2(N__32535),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_11_27_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_11_27_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_11_27_6  (
            .in0(_gnd_net_),
            .in1(N__32523),
            .in2(N__32514),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_11_27_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_11_27_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_11_27_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_11_27_7  (
            .in0(_gnd_net_),
            .in1(N__32628),
            .in2(N__32550),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_28_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_28_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_11_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32517),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_11_28_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_11_28_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_11_28_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_11_28_2  (
            .in0(_gnd_net_),
            .in1(N__36966),
            .in2(_gnd_net_),
            .in3(N__36896),
            .lcout(\phase_controller_inst1.stoper_tr.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_28_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_28_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_28_3 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_11_28_3  (
            .in0(N__34944),
            .in1(N__35786),
            .in2(_gnd_net_),
            .in3(N__35814),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_28_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_28_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_28_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_28_5  (
            .in0(N__33776),
            .in1(N__35938),
            .in2(N__35042),
            .in3(N__35485),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_28_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_28_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_28_6 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_28_6  (
            .in0(N__35114),
            .in1(N__35007),
            .in2(N__35511),
            .in3(N__35531),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_28_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_28_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_28_7 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_28_7  (
            .in0(N__33777),
            .in1(N__35939),
            .in2(N__35043),
            .in3(N__35486),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_29_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_29_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_29_0 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_29_0  (
            .in0(N__35006),
            .in1(N__35506),
            .in2(N__35115),
            .in3(N__35530),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_11_29_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_11_29_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_11_29_2 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_11_29_2  (
            .in0(N__35896),
            .in1(N__35132),
            .in2(N__34971),
            .in3(N__35920),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_29_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_29_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_29_7 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_11_29_7  (
            .in0(N__35756),
            .in1(N__35597),
            .in2(_gnd_net_),
            .in3(N__34945),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_30_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_30_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_30_3 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_11_30_3  (
            .in0(N__35133),
            .in1(N__34970),
            .in2(N__35901),
            .in3(N__35921),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_30_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_30_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_30_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_30_6  (
            .in0(N__41171),
            .in1(N__40893),
            .in2(_gnd_net_),
            .in3(N__40925),
            .lcout(\current_shift_inst.timer_s1.N_154_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_11_30_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_11_30_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_11_30_7 .LUT_INIT=16'b1111000011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_11_30_7  (
            .in0(_gnd_net_),
            .in1(N__35755),
            .in2(N__34949),
            .in3(N__35596),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_6_2 .LUT_INIT=16'b1100110000001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__32799),
            .in2(N__38212),
            .in3(N__32815),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_12_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_12_6_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_12_6_4  (
            .in0(N__52082),
            .in1(N__32798),
            .in2(_gnd_net_),
            .in3(N__38214),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_12_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_12_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_3_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37293),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52460),
            .ce(N__36314),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_12_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_12_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_5_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37233),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52460),
            .ce(N__36314),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_12_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_12_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_2_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37323),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52460),
            .ce(N__36314),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_12_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_12_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_1_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37353),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52460),
            .ce(N__36314),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_12_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_12_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_8_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37152),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52456),
            .ce(N__36324),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_12_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_12_9_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_12_9_0  (
            .in0(N__36462),
            .in1(N__32715),
            .in2(N__36360),
            .in3(N__32697),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_12_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_12_9_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_12_9_2  (
            .in0(N__36461),
            .in1(N__32714),
            .in2(N__36359),
            .in3(N__32696),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_12_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_12_9_4 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_12_9_4  (
            .in0(N__32972),
            .in1(N__36042),
            .in2(N__36447),
            .in3(N__32954),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_12_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_12_9_6 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_12_9_6  (
            .in0(N__32971),
            .in1(N__36041),
            .in2(N__36446),
            .in3(N__32953),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_10_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_10_0  (
            .in0(N__36098),
            .in1(N__36248),
            .in2(_gnd_net_),
            .in3(N__38914),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_10_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_10_2  (
            .in0(N__36097),
            .in1(N__36247),
            .in2(_gnd_net_),
            .in3(N__38913),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_12_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_4_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37263),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52437),
            .ce(N__36332),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_12_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_9_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37548),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52437),
            .ce(N__36332),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_12_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_13_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37461),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52437),
            .ce(N__36332),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_12_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_12_11_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_17_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__37377),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52437),
            .ce(N__36332),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_12_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_12_12_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_25_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__37569),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52432),
            .ce(N__36333),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_12_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_12_12_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_12_12_4  (
            .in0(N__32877),
            .in1(N__36029),
            .in2(N__32850),
            .in3(N__36476),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_12_13_2  (
            .in0(N__33100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52427),
            .ce(),
            .sr(N__51953));
    defparam \phase_controller_inst1.state_1_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_13_3 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_13_3  (
            .in0(N__37072),
            .in1(N__38246),
            .in2(N__36758),
            .in3(N__36787),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52427),
            .ce(),
            .sr(N__51953));
    defparam \phase_controller_inst1.start_timer_hc_LC_12_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_13_6 .LUT_INIT=16'b1010101011111000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_12_13_6  (
            .in0(N__41217),
            .in1(N__36646),
            .in2(N__33104),
            .in3(N__36753),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52427),
            .ce(),
            .sr(N__51953));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_12_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_10_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37524),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_12_14_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_0_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__42297),
            .in2(_gnd_net_),
            .in3(N__39615),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_12_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_11_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37503),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_12_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_12_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_24_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37590),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_12_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_12_14_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_6_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__37202),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_12_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_12_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37482),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_12_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_12_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_14_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37440),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52421),
            .ce(N__36334),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36844),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33468),
            .ce(),
            .sr(N__51962));
    defparam \delay_measurement_inst.start_timer_tr_LC_12_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_12_15_5  (
            .in0(N__36845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33468),
            .ce(),
            .sr(N__51962));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_16_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__33136),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__37737),
            .in2(_gnd_net_),
            .in3(N__36817),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_157_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_16_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_12_16_2  (
            .in0(N__34855),
            .in1(N__34209),
            .in2(N__33453),
            .in3(N__33410),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_16_5 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_12_16_5  (
            .in0(N__34211),
            .in1(N__33374),
            .in2(N__33332),
            .in3(N__34857),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_12_16_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_12_16_7  (
            .in0(N__34210),
            .in1(N__34856),
            .in2(N__33281),
            .in3(N__33248),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33189),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52406),
            .ce(N__33757),
            .sr(N__51972));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_17_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_17_5  (
            .in0(N__34208),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33722),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33915),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_18_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_12_18_5  (
            .in0(N__34244),
            .in1(N__34858),
            .in2(N__33689),
            .in3(N__33638),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__36759),
            .in2(_gnd_net_),
            .in3(N__36794),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_12_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_12_19_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_12_19_2  (
            .in0(N__52085),
            .in1(N__37013),
            .in2(_gnd_net_),
            .in3(N__36974),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_12_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_12_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__42503),
            .in2(_gnd_net_),
            .in3(N__42522),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33588),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_12_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_12_19_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_12_19_5  (
            .in0(N__34907),
            .in1(N__34246),
            .in2(N__33549),
            .in3(N__33509),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_12_19_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_12_19_7  (
            .in0(N__34906),
            .in1(N__34245),
            .in2(N__33921),
            .in3(N__33882),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37412),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52391),
            .ce(N__38374),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37517),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52391),
            .ce(N__38374),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37475),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52391),
            .ce(N__38374),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_12_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_12_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_7_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37172),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_12_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_16_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37391),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37496),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37433),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_12_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_12_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_22_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37625),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_12_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_12_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_13_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37454),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_12_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_12_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_23_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37604),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52388),
            .ce(N__38405),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_12_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_12_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_27_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37757),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52383),
            .ce(N__38423),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_22_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37541),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52383),
            .ce(N__38423),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_12_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_12_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_18_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37694),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52383),
            .ce(N__38423),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_12_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_12_22_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_12_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_21_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37646),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52383),
            .ce(N__38423),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_12_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_12_23_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_0_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__42296),
            .in2(_gnd_net_),
            .in3(N__39614),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52380),
            .ce(N__38409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_12_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_12_23_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_12_23_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_25_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__37562),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52380),
            .ce(N__38409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40463),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52380),
            .ce(N__38409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_12_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_12_23_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_17_LC_12_23_4  (
            .in0(N__37373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52380),
            .ce(N__38409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_12_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_12_23_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_12_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_26_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37778),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52380),
            .ce(N__38409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_12_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_12_23_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_24_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__37583),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52380),
            .ce(N__38409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_12_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_12_24_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_12_24_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_20_LC_12_24_0  (
            .in0(N__37676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52376),
            .ce(N__38404),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_12_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_12_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_5_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37229),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52376),
            .ce(N__38404),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_12_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_12_24_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_12_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_3_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37289),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52376),
            .ce(N__38404),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_12_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_12_25_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_12_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37352),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52373),
            .ce(N__38419),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_12_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_12_25_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_12_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_2_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37319),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52373),
            .ce(N__38419),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_12_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_12_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_6_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37203),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52373),
            .ce(N__38419),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_25_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37148),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52373),
            .ce(N__38419),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_12_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_12_25_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_12_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_4_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37262),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52373),
            .ce(N__38419),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_12_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_12_26_2 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_12_26_2  (
            .in0(N__35840),
            .in1(N__35301),
            .in2(N__35877),
            .in3(N__35285),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_12_27_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_12_27_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_12_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_0_LC_12_27_0  (
            .in0(N__35705),
            .in1(N__35246),
            .in2(N__35262),
            .in3(N__35261),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_27_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_0 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_12_27_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_12_27_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_12_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_1_LC_12_27_1  (
            .in0(N__35733),
            .in1(N__35231),
            .in2(_gnd_net_),
            .in3(N__35217),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_1 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_12_27_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_12_27_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_12_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_2_LC_12_27_2  (
            .in0(N__35706),
            .in1(N__35210),
            .in2(_gnd_net_),
            .in3(N__35196),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_2 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_12_27_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_12_27_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_12_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_3_LC_12_27_3  (
            .in0(N__35734),
            .in1(N__35189),
            .in2(_gnd_net_),
            .in3(N__35175),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_3 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_12_27_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_12_27_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_12_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_4_LC_12_27_4  (
            .in0(N__35707),
            .in1(N__35171),
            .in2(_gnd_net_),
            .in3(N__35157),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_4 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_12_27_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_12_27_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_12_27_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_5_LC_12_27_5  (
            .in0(N__35735),
            .in1(N__35150),
            .in2(_gnd_net_),
            .in3(N__35136),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_5 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_12_27_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_12_27_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_12_27_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_6_LC_12_27_6  (
            .in0(N__35708),
            .in1(N__35468),
            .in2(_gnd_net_),
            .in3(N__35454),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_6 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_12_27_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_12_27_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_12_27_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_7_LC_12_27_7  (
            .in0(N__35736),
            .in1(N__35450),
            .in2(_gnd_net_),
            .in3(N__35436),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_7 ),
            .clk(N__52370),
            .ce(N__35580),
            .sr(N__52034));
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_12_28_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_12_28_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_12_28_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_8_LC_12_28_0  (
            .in0(N__35712),
            .in1(N__35432),
            .in2(_gnd_net_),
            .in3(N__35418),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_28_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_8 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_12_28_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_12_28_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_12_28_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_9_LC_12_28_1  (
            .in0(N__35729),
            .in1(N__35414),
            .in2(_gnd_net_),
            .in3(N__35400),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_9 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_12_28_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_12_28_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_12_28_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_10_LC_12_28_2  (
            .in0(N__35709),
            .in1(N__35396),
            .in2(_gnd_net_),
            .in3(N__35382),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_10 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_12_28_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_12_28_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_12_28_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_11_LC_12_28_3  (
            .in0(N__35726),
            .in1(N__35378),
            .in2(_gnd_net_),
            .in3(N__35364),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_11 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_12_28_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_12_28_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_12_28_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_12_LC_12_28_4  (
            .in0(N__35710),
            .in1(N__35360),
            .in2(_gnd_net_),
            .in3(N__35346),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_12 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_12_28_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_12_28_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_12_28_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_13_LC_12_28_5  (
            .in0(N__35727),
            .in1(N__35342),
            .in2(_gnd_net_),
            .in3(N__35328),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_13 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_12_28_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_12_28_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_12_28_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_14_LC_12_28_6  (
            .in0(N__35711),
            .in1(N__35324),
            .in2(_gnd_net_),
            .in3(N__35310),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_14 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_12_28_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_12_28_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_12_28_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_15_LC_12_28_7  (
            .in0(N__35728),
            .in1(N__35561),
            .in2(_gnd_net_),
            .in3(N__35547),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_15 ),
            .clk(N__52367),
            .ce(N__35579),
            .sr(N__52038));
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_12_29_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_12_29_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_12_29_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_16_LC_12_29_0  (
            .in0(N__35713),
            .in1(N__37867),
            .in2(_gnd_net_),
            .in3(N__35544),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_29_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_16 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_12_29_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_12_29_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_12_29_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_17_LC_12_29_1  (
            .in0(N__35717),
            .in1(N__37921),
            .in2(_gnd_net_),
            .in3(N__35541),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_17 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_12_29_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_12_29_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_12_29_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_18_LC_12_29_2  (
            .in0(N__35714),
            .in1(N__38343),
            .in2(_gnd_net_),
            .in3(N__35538),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_18 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_12_29_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_12_29_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_12_29_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_19_LC_12_29_3  (
            .in0(N__35718),
            .in1(N__38300),
            .in2(_gnd_net_),
            .in3(N__35535),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_19 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_12_29_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_12_29_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_12_29_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_20_LC_12_29_4  (
            .in0(N__35715),
            .in1(N__35532),
            .in2(_gnd_net_),
            .in3(N__35514),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_20 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_12_29_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_12_29_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_12_29_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_21_LC_12_29_5  (
            .in0(N__35719),
            .in1(N__35510),
            .in2(_gnd_net_),
            .in3(N__35490),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_21 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_12_29_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_12_29_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_12_29_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_22_LC_12_29_6  (
            .in0(N__35716),
            .in1(N__35487),
            .in2(_gnd_net_),
            .in3(N__35472),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_22 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_12_29_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_12_29_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_12_29_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_23_LC_12_29_7  (
            .in0(N__35720),
            .in1(N__35940),
            .in2(_gnd_net_),
            .in3(N__35925),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_23 ),
            .clk(N__52366),
            .ce(N__35578),
            .sr(N__52043));
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_12_30_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_12_30_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_12_30_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_24_LC_12_30_0  (
            .in0(N__35721),
            .in1(N__35922),
            .in2(_gnd_net_),
            .in3(N__35904),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_12_30_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_24 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_12_30_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_12_30_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_12_30_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_25_LC_12_30_1  (
            .in0(N__35730),
            .in1(N__35900),
            .in2(_gnd_net_),
            .in3(N__35880),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_25 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_12_30_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_12_30_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_12_30_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_26_LC_12_30_2  (
            .in0(N__35722),
            .in1(N__35863),
            .in2(_gnd_net_),
            .in3(N__35847),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_26 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_12_30_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_12_30_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_12_30_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_27_LC_12_30_3  (
            .in0(N__35731),
            .in1(N__35839),
            .in2(_gnd_net_),
            .in3(N__35817),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_27 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_12_30_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_12_30_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_12_30_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_28_LC_12_30_4  (
            .in0(N__35723),
            .in1(N__35806),
            .in2(_gnd_net_),
            .in3(N__35790),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_28 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_12_30_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_12_30_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_12_30_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_29_LC_12_30_5  (
            .in0(N__35732),
            .in1(N__35782),
            .in2(_gnd_net_),
            .in3(N__35760),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_29 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_12_30_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_12_30_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_12_30_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_30_LC_12_30_6  (
            .in0(N__35724),
            .in1(N__35757),
            .in2(_gnd_net_),
            .in3(N__35739),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_30 ),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_12_30_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_12_30_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_12_30_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_31_LC_12_30_7  (
            .in0(N__35598),
            .in1(N__35725),
            .in2(_gnd_net_),
            .in3(N__35601),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52365),
            .ce(N__35577),
            .sr(N__52045));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_13_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_13_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38213),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_13_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_13_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_0_LC_13_7_0  (
            .in0(N__36193),
            .in1(N__38151),
            .in2(N__38169),
            .in3(N__38165),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_0 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_13_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_13_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_1_LC_13_7_1  (
            .in0(N__36225),
            .in1(N__38133),
            .in2(_gnd_net_),
            .in3(N__35961),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_1 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_13_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_13_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_2_LC_13_7_2  (
            .in0(N__36194),
            .in1(N__38604),
            .in2(_gnd_net_),
            .in3(N__35958),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_2 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_13_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_13_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_3_LC_13_7_3  (
            .in0(N__36226),
            .in1(N__38586),
            .in2(_gnd_net_),
            .in3(N__35955),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_3 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_13_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_13_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_4_LC_13_7_4  (
            .in0(N__36195),
            .in1(N__38568),
            .in2(_gnd_net_),
            .in3(N__35952),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_4 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_13_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_13_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_5_LC_13_7_5  (
            .in0(N__36227),
            .in1(N__38550),
            .in2(_gnd_net_),
            .in3(N__35949),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_5 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_13_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_13_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_6_LC_13_7_6  (
            .in0(N__36196),
            .in1(N__38529),
            .in2(_gnd_net_),
            .in3(N__35946),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_6 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_13_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_13_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_7_LC_13_7_7  (
            .in0(N__36228),
            .in1(N__38505),
            .in2(_gnd_net_),
            .in3(N__35943),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_7 ),
            .clk(N__52467),
            .ce(N__36058),
            .sr(N__51928));
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_13_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_13_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_8_LC_13_8_0  (
            .in0(N__36205),
            .in1(N__38484),
            .in2(_gnd_net_),
            .in3(N__35988),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_8 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_13_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_13_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_9_LC_13_8_1  (
            .in0(N__36224),
            .in1(N__38463),
            .in2(_gnd_net_),
            .in3(N__35985),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_9 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_13_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_13_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_10_LC_13_8_2  (
            .in0(N__36202),
            .in1(N__38733),
            .in2(_gnd_net_),
            .in3(N__35982),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_10 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_13_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_13_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_11_LC_13_8_3  (
            .in0(N__36221),
            .in1(N__38712),
            .in2(_gnd_net_),
            .in3(N__35979),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_11 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_13_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_13_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_12_LC_13_8_4  (
            .in0(N__36203),
            .in1(N__38691),
            .in2(_gnd_net_),
            .in3(N__35976),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_12 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_13_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_13_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_13_LC_13_8_5  (
            .in0(N__36222),
            .in1(N__38667),
            .in2(_gnd_net_),
            .in3(N__35973),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_13 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_13_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_13_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_14_LC_13_8_6  (
            .in0(N__36204),
            .in1(N__38646),
            .in2(_gnd_net_),
            .in3(N__35970),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_14 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_13_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_13_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_15_LC_13_8_7  (
            .in0(N__36223),
            .in1(N__38625),
            .in2(_gnd_net_),
            .in3(N__35967),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_15 ),
            .clk(N__52462),
            .ce(N__36076),
            .sr(N__51933));
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_13_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_13_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_16_LC_13_9_0  (
            .in0(N__36206),
            .in1(N__49957),
            .in2(_gnd_net_),
            .in3(N__35964),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_16 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_13_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_13_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_17_LC_13_9_1  (
            .in0(N__36210),
            .in1(N__49981),
            .in2(_gnd_net_),
            .in3(N__36015),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_17 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_13_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_13_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_18_LC_13_9_2  (
            .in0(N__36207),
            .in1(N__49843),
            .in2(_gnd_net_),
            .in3(N__36012),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_18 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_13_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_13_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_19_LC_13_9_3  (
            .in0(N__36211),
            .in1(N__49865),
            .in2(_gnd_net_),
            .in3(N__36009),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_19 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_13_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_13_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_20_LC_13_9_4  (
            .in0(N__36208),
            .in1(N__41288),
            .in2(_gnd_net_),
            .in3(N__36006),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_20 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_13_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_13_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_21_LC_13_9_5  (
            .in0(N__36212),
            .in1(N__41315),
            .in2(_gnd_net_),
            .in3(N__36003),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_21 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_13_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_13_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_22_LC_13_9_6  (
            .in0(N__36209),
            .in1(N__41642),
            .in2(_gnd_net_),
            .in3(N__36000),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_22 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_13_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_13_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_23_LC_13_9_7  (
            .in0(N__36213),
            .in1(N__41678),
            .in2(_gnd_net_),
            .in3(N__35997),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_23 ),
            .clk(N__52458),
            .ce(N__36077),
            .sr(N__51934));
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_13_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_13_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_24_LC_13_10_0  (
            .in0(N__36197),
            .in1(N__49771),
            .in2(_gnd_net_),
            .in3(N__35994),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_24 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_13_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_13_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_25_LC_13_10_1  (
            .in0(N__36229),
            .in1(N__49789),
            .in2(_gnd_net_),
            .in3(N__35991),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_25 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_13_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_13_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_26_LC_13_10_2  (
            .in0(N__36198),
            .in1(N__50305),
            .in2(_gnd_net_),
            .in3(N__36261),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_26 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_13_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_13_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_27_LC_13_10_3  (
            .in0(N__36230),
            .in1(N__50276),
            .in2(_gnd_net_),
            .in3(N__36258),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_27 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_13_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_13_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_28_LC_13_10_4  (
            .in0(N__36199),
            .in1(N__38934),
            .in2(_gnd_net_),
            .in3(N__36255),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_28 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_13_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_13_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_29_LC_13_10_5  (
            .in0(N__36231),
            .in1(N__38898),
            .in2(_gnd_net_),
            .in3(N__36252),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_29 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_13_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_13_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_30_LC_13_10_6  (
            .in0(N__36200),
            .in1(N__36249),
            .in2(_gnd_net_),
            .in3(N__36234),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_29 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_30 ),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_13_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_13_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_13_10_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_31_LC_13_10_7  (
            .in0(N__36099),
            .in1(N__36201),
            .in2(_gnd_net_),
            .in3(N__36102),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52452),
            .ce(N__36084),
            .sr(N__51940));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_13_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_13_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_28_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47667),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52445),
            .ce(N__50155),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_13_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_22_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37632),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52439),
            .ce(N__36335),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_13_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_26_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37785),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52439),
            .ce(N__36335),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_13_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_13_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_15_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37419),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52439),
            .ce(N__36335),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_13_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_27_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37764),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52439),
            .ce(N__36335),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_13_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_20_LC_13_12_7  (
            .in0(N__37677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52439),
            .ce(N__36335),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_13_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_13_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_23_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37611),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52434),
            .ce(N__36339),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_13_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_7_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37176),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52434),
            .ce(N__36339),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_13_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_18_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37698),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52434),
            .ce(N__36339),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_13_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_16_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37398),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52434),
            .ce(N__36339),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_13_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_13_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_19_LC_13_13_5  (
            .in0(N__38442),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52434),
            .ce(N__36339),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_13_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_13_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_21_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37653),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52434),
            .ce(N__36339),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_13_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_13_14_1 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_13_14_1  (
            .in0(N__36653),
            .in1(N__36754),
            .in2(N__41218),
            .in3(N__36795),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52429),
            .ce(),
            .sr(N__51954));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_13_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_13_14_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_13_14_5  (
            .in0(N__39157),
            .in1(N__39881),
            .in2(_gnd_net_),
            .in3(N__39909),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_13_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_13_14_6 .LUT_INIT=16'b1100110111001101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_13_14_6  (
            .in0(N__39908),
            .in1(N__39156),
            .in2(N__39885),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_13_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_13_15_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_13_15_0  (
            .in0(N__39704),
            .in1(N__39857),
            .in2(_gnd_net_),
            .in3(N__39158),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47660),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52422),
            .ce(N__43467),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_16_1 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_13_16_1  (
            .in0(N__37738),
            .in1(N__36843),
            .in2(_gnd_net_),
            .in3(N__36821),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52417),
            .ce(),
            .sr(N__51963));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_16_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__36728),
            .in2(_gnd_net_),
            .in3(N__36707),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52417),
            .ce(),
            .sr(N__51963));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_17_0 .LUT_INIT=16'b0100010111001111;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_13_17_0  (
            .in0(N__37102),
            .in1(N__36657),
            .in2(N__41211),
            .in3(N__37091),
            .lcout(),
            .ltout(\phase_controller_inst1.state_ns_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_13_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_17_1 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_17_1  (
            .in0(N__36604),
            .in1(N__36534),
            .in2(N__36516),
            .in3(N__36513),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52411),
            .ce(),
            .sr(N__51966));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_17_3 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_17_3  (
            .in0(N__37122),
            .in1(N__37106),
            .in2(N__36881),
            .in3(N__36911),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52411),
            .ce(),
            .sr(N__51966));
    defparam \phase_controller_inst1.state_0_LC_13_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_13_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_13_17_4 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_inst1.state_0_LC_13_17_4  (
            .in0(N__37082),
            .in1(N__38260),
            .in2(N__37107),
            .in3(N__37092),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52411),
            .ce(),
            .sr(N__51966));
    defparam \phase_controller_inst1.start_timer_tr_LC_13_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_17_5 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_13_17_5  (
            .in0(N__38261),
            .in1(N__37032),
            .in2(N__37083),
            .in3(N__37047),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52411),
            .ce(),
            .sr(N__51966));
    defparam \phase_controller_inst1.stoper_tr.running_LC_13_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_13_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_13_17_7 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_13_17_7  (
            .in0(N__36877),
            .in1(N__37031),
            .in2(N__36978),
            .in3(N__36912),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52411),
            .ce(),
            .sr(N__51966));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_13_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_13_18_2  (
            .in0(N__44154),
            .in1(N__43953),
            .in2(N__44205),
            .in3(N__43932),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_13_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_13_18_3  (
            .in0(N__44177),
            .in1(N__44228),
            .in2(N__36858),
            .in3(N__36855),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_18_4 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_18_4  (
            .in0(N__37740),
            .in1(_gnd_net_),
            .in2(N__36849),
            .in3(N__36822),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_158_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_18_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__39210),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_13_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_13_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__36801),
            .in2(N__39604),
            .in3(N__42295),
            .lcout(\phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_13_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_13_19_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_13_19_1  (
            .in0(N__39579),
            .in1(N__39578),
            .in2(N__46684),
            .in3(N__37326),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_1),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_13_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_13_19_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_13_19_2  (
            .in0(N__40050),
            .in1(N__40049),
            .in2(N__46688),
            .in3(N__37296),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_2),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_13_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_13_19_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_13_19_3  (
            .in0(N__40035),
            .in1(N__40034),
            .in2(N__46685),
            .in3(N__37266),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_3),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_13_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_13_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_13_19_4  (
            .in0(N__40020),
            .in1(N__40019),
            .in2(N__46689),
            .in3(N__37236),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_4),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_13_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_13_19_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_13_19_5  (
            .in0(N__40005),
            .in1(N__40004),
            .in2(N__46686),
            .in3(N__37206),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_5),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_13_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_13_19_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_13_19_6  (
            .in0(N__39978),
            .in1(N__39977),
            .in2(N__46690),
            .in3(N__37179),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_6),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_13_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_13_19_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_13_19_7  (
            .in0(N__39957),
            .in1(N__39956),
            .in2(N__46687),
            .in3(N__37155),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_7),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_13_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_13_20_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_13_20_0  (
            .in0(N__39939),
            .in1(N__39938),
            .in2(N__46842),
            .in3(N__37125),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_8),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_13_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_13_20_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_13_20_1  (
            .in0(N__39924),
            .in1(N__39923),
            .in2(N__46839),
            .in3(N__37527),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_9),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_13_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_13_20_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_13_20_2  (
            .in0(N__40200),
            .in1(N__40199),
            .in2(N__46843),
            .in3(N__37506),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_10),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_13_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_13_20_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_13_20_3  (
            .in0(N__40185),
            .in1(N__40184),
            .in2(N__46836),
            .in3(N__37485),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_11),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_13_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_13_20_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_13_20_4  (
            .in0(N__40170),
            .in1(N__40169),
            .in2(N__46840),
            .in3(N__37464),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_12),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_13_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_13_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_13_20_5  (
            .in0(N__40155),
            .in1(N__40154),
            .in2(N__46837),
            .in3(N__37443),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_13),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_13_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_13_20_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_13_20_6  (
            .in0(N__40140),
            .in1(N__40139),
            .in2(N__46841),
            .in3(N__37422),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_14),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_13_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_13_20_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_13_20_7  (
            .in0(N__40119),
            .in1(N__40118),
            .in2(N__46838),
            .in3(N__37401),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_15),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_13_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_13_21_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_13_21_0  (
            .in0(N__40101),
            .in1(N__40100),
            .in2(N__46844),
            .in3(N__37380),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_16),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_13_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_13_21_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_13_21_1  (
            .in0(N__40082),
            .in1(N__40086),
            .in2(N__46872),
            .in3(N__37356),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_17),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_13_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_13_21_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_13_21_2  (
            .in0(N__40065),
            .in1(N__40064),
            .in2(N__46845),
            .in3(N__37683),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_18),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_13_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_13_21_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_13_21_3  (
            .in0(N__40329),
            .in1(N__40328),
            .in2(N__46873),
            .in3(N__37680),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_19),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_13_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_13_21_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_13_21_4  (
            .in0(N__40314),
            .in1(N__40313),
            .in2(N__46846),
            .in3(N__37656),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_20),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_13_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_13_21_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_13_21_5  (
            .in0(N__40299),
            .in1(N__40298),
            .in2(N__46874),
            .in3(N__37635),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_21),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_13_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_13_21_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_13_21_6  (
            .in0(N__40284),
            .in1(N__40283),
            .in2(N__46847),
            .in3(N__37614),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_22),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_13_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_13_21_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_13_21_7  (
            .in0(N__40263),
            .in1(N__40262),
            .in2(N__46875),
            .in3(N__37593),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_23),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_13_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_13_22_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_13_22_0  (
            .in0(N__40245),
            .in1(N__40244),
            .in2(N__46876),
            .in3(N__37572),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_24),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_13_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_13_22_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_13_22_1  (
            .in0(N__40230),
            .in1(N__40229),
            .in2(N__46878),
            .in3(N__37551),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_25),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_13_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_13_22_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_13_22_2  (
            .in0(N__40215),
            .in1(N__40214),
            .in2(N__46877),
            .in3(N__37767),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_26),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_13_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_13_22_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_13_22_3  (
            .in0(N__40494),
            .in1(N__40493),
            .in2(N__46879),
            .in3(N__37746),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_27),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_13_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37743),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37739),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_23_0  (
            .in0(N__38054),
            .in1(N__42223),
            .in2(_gnd_net_),
            .in3(N__37713),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_23_1  (
            .in0(N__38088),
            .in1(N__42175),
            .in2(_gnd_net_),
            .in3(N__37710),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_23_2  (
            .in0(N__38055),
            .in1(N__40443),
            .in2(_gnd_net_),
            .in3(N__37707),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_23_3  (
            .in0(N__38089),
            .in1(N__40421),
            .in2(_gnd_net_),
            .in3(N__37704),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_23_4  (
            .in0(N__38056),
            .in1(N__40399),
            .in2(_gnd_net_),
            .in3(N__37701),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_23_5  (
            .in0(N__38090),
            .in1(N__40373),
            .in2(_gnd_net_),
            .in3(N__37812),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_23_6  (
            .in0(N__38057),
            .in1(N__40349),
            .in2(_gnd_net_),
            .in3(N__37809),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_23_7  (
            .in0(N__38091),
            .in1(N__40679),
            .in2(_gnd_net_),
            .in3(N__37806),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__52385),
            .ce(N__37972),
            .sr(N__51999));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_24_0  (
            .in0(N__38075),
            .in1(N__40655),
            .in2(_gnd_net_),
            .in3(N__37803),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_24_1  (
            .in0(N__38087),
            .in1(N__40634),
            .in2(_gnd_net_),
            .in3(N__37800),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_24_2  (
            .in0(N__38072),
            .in1(N__40610),
            .in2(_gnd_net_),
            .in3(N__37797),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_24_3  (
            .in0(N__38084),
            .in1(N__40588),
            .in2(_gnd_net_),
            .in3(N__37794),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_24_4  (
            .in0(N__38073),
            .in1(N__40562),
            .in2(_gnd_net_),
            .in3(N__37791),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_24_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_24_5  (
            .in0(N__38085),
            .in1(N__40538),
            .in2(_gnd_net_),
            .in3(N__37788),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_24_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_24_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_24_6  (
            .in0(N__38074),
            .in1(N__40514),
            .in2(_gnd_net_),
            .in3(N__37839),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_24_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_24_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_24_7  (
            .in0(N__38086),
            .in1(N__40865),
            .in2(_gnd_net_),
            .in3(N__37836),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__52381),
            .ce(N__37968),
            .sr(N__52005));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_25_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_25_0  (
            .in0(N__38076),
            .in1(N__40841),
            .in2(_gnd_net_),
            .in3(N__37833),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_25_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_25_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_25_1  (
            .in0(N__38080),
            .in1(N__40817),
            .in2(_gnd_net_),
            .in3(N__37830),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_25_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_25_2  (
            .in0(N__38077),
            .in1(N__40797),
            .in2(_gnd_net_),
            .in3(N__37827),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_25_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_25_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_25_3  (
            .in0(N__38081),
            .in1(N__40775),
            .in2(_gnd_net_),
            .in3(N__37824),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_25_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_25_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_25_4  (
            .in0(N__38078),
            .in1(N__40753),
            .in2(_gnd_net_),
            .in3(N__37821),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_25_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_25_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_25_5  (
            .in0(N__38082),
            .in1(N__40727),
            .in2(_gnd_net_),
            .in3(N__37818),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_25_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_25_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_25_6  (
            .in0(N__38079),
            .in1(N__40703),
            .in2(_gnd_net_),
            .in3(N__37815),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_25_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_25_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_25_7  (
            .in0(N__38083),
            .in1(N__41069),
            .in2(_gnd_net_),
            .in3(N__38115),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__52377),
            .ce(N__37973),
            .sr(N__52012));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_26_0  (
            .in0(N__38092),
            .in1(N__41045),
            .in2(_gnd_net_),
            .in3(N__38112),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__52374),
            .ce(N__37974),
            .sr(N__52021));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_26_1  (
            .in0(N__38096),
            .in1(N__41024),
            .in2(_gnd_net_),
            .in3(N__38109),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__52374),
            .ce(N__37974),
            .sr(N__52021));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_26_2  (
            .in0(N__38093),
            .in1(N__40988),
            .in2(_gnd_net_),
            .in3(N__38106),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__52374),
            .ce(N__37974),
            .sr(N__52021));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_26_3  (
            .in0(N__38097),
            .in1(N__40954),
            .in2(_gnd_net_),
            .in3(N__38103),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__52374),
            .ce(N__37974),
            .sr(N__52021));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_26_4  (
            .in0(N__38094),
            .in1(N__41004),
            .in2(_gnd_net_),
            .in3(N__38100),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__52374),
            .ce(N__37974),
            .sr(N__52021));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_26_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_26_5  (
            .in0(N__40968),
            .in1(N__38095),
            .in2(_gnd_net_),
            .in3(N__37977),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52374),
            .ce(N__37974),
            .sr(N__52021));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_13_27_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_13_27_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_13_27_0  (
            .in0(N__37923),
            .in1(N__37905),
            .in2(N__37890),
            .in3(N__37869),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_13_27_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_13_27_2 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_13_27_2  (
            .in0(N__37922),
            .in1(N__37904),
            .in2(N__37889),
            .in3(N__37868),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_13_27_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_13_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_19_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38441),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52372),
            .ce(N__38424),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_13_28_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_13_28_2 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_13_28_2  (
            .in0(N__38327),
            .in1(N__38312),
            .in2(N__38301),
            .in3(N__38341),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_13_28_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_13_28_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_13_28_3 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_13_28_3  (
            .in0(N__38342),
            .in1(N__38328),
            .in2(N__38313),
            .in3(N__38299),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_29_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_29_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_29_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_29_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38271),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52368),
            .ce(),
            .sr(N__52039));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_30_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_30_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_30_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_30_0  (
            .in0(_gnd_net_),
            .in1(N__40914),
            .in2(_gnd_net_),
            .in3(N__40887),
            .lcout(\current_shift_inst.timer_s1.N_153_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_14_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_14_7_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__38219),
            .in2(_gnd_net_),
            .in3(N__38762),
            .lcout(\phase_controller_inst2.stoper_hc.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_14_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_14_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__38139),
            .in2(N__41148),
            .in3(N__38150),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_0 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_14_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_14_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__38121),
            .in2(N__41121),
            .in3(N__38132),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_14_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_14_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__38592),
            .in2(N__41112),
            .in3(N__38603),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_14_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_14_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__38574),
            .in2(N__41139),
            .in3(N__38585),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_14_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_14_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__38556),
            .in2(N__41130),
            .in3(N__38567),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_14_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_14_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__43245),
            .in2(N__38538),
            .in3(N__38549),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_14_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_14_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__41103),
            .in2(N__38517),
            .in3(N__38528),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_14_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_14_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__43236),
            .in2(N__38493),
            .in3(N__38504),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_14_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_14_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__43383),
            .in2(N__38472),
            .in3(N__38483),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_8 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_14_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_14_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__43200),
            .in2(N__38451),
            .in3(N__38462),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_14_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_14_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__43227),
            .in2(N__38721),
            .in3(N__38732),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_14_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_14_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__43269),
            .in2(N__38700),
            .in3(N__38711),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_14_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_14_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_14_9_4  (
            .in0(N__38690),
            .in1(N__43209),
            .in2(N__38679),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_14_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_14_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__43392),
            .in2(N__38655),
            .in3(N__38666),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_14_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_14_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__43257),
            .in2(N__38634),
            .in3(N__38645),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_14_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_14_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__43218),
            .in2(N__38613),
            .in3(N__38624),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_14_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_14_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__50004),
            .in2(N__49938),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_14_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_14_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__49818),
            .in2(N__49896),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_14_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_14_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__41274),
            .in2(N__41343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_14_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_14_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__41259),
            .in2(N__41628),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_14_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_14_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(N__49755),
            .in2(N__49806),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_14_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_14_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__49746),
            .in2(N__50262),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_14_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_14_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__38883),
            .in2(N__38745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_14_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_14_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__38796),
            .in2(N__38787),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38775),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_14_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_14_11_1 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_14_11_1  (
            .in0(N__38896),
            .in1(N__38918),
            .in2(_gnd_net_),
            .in3(N__38932),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_11_2 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_11_2  (
            .in0(N__41612),
            .in1(N__43500),
            .in2(N__41583),
            .in3(N__43485),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_14_11_6 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_14_11_6  (
            .in0(N__38933),
            .in1(_gnd_net_),
            .in2(N__38919),
            .in3(N__38897),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_12_0  (
            .in0(N__39087),
            .in1(N__38877),
            .in2(N__38862),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_0 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__41373),
            .in2(N__38853),
            .in3(N__39072),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__41352),
            .in2(N__38844),
            .in3(N__39378),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__43374),
            .in2(N__38835),
            .in3(N__39360),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__43551),
            .in2(N__38826),
            .in3(N__39342),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_12_5  (
            .in0(N__39324),
            .in1(N__43350),
            .in2(N__38814),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_12_6  (
            .in0(N__39306),
            .in1(N__41097),
            .in2(N__38805),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_12_7  (
            .in0(N__39288),
            .in1(N__43515),
            .in2(N__39012),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__41085),
            .in2(N__39003),
            .in3(N__39270),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_8 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__43296),
            .in2(N__38994),
            .in3(N__39252),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__43284),
            .in2(N__38985),
            .in3(N__39498),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__41364),
            .in2(N__38976),
            .in3(N__39480),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_13_4  (
            .in0(N__39462),
            .in1(N__41385),
            .in2(N__38964),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_13_5  (
            .in0(N__39441),
            .in1(N__43338),
            .in2(N__38952),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_13_6  (
            .in0(N__39423),
            .in1(N__43326),
            .in2(N__38943),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_13_7  (
            .in0(N__39405),
            .in1(N__43362),
            .in2(N__39054),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__41838),
            .in2(N__41784),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__41766),
            .in2(N__41703),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__41535),
            .in2(N__41466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__41454),
            .in2(N__41859),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__39045),
            .in2(N__41550),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__39120),
            .in2(N__39129),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__39036),
            .in2(N__39030),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__39018),
            .in2(N__39138),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39234),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ),
            .ltout(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_15_1 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39213),
            .in3(N__39208),
            .lcout(\phase_controller_inst1.stoper_hc.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_14_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_14_15_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_14_15_3  (
            .in0(N__39705),
            .in1(N__39858),
            .in2(_gnd_net_),
            .in3(N__39159),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_15_4 .LUT_INIT=16'b0100000011011100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_15_4  (
            .in0(N__39543),
            .in1(N__43313),
            .in2(N__43578),
            .in3(N__39522),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_15_5 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_15_5  (
            .in0(N__39521),
            .in1(N__43574),
            .in2(N__43314),
            .in3(N__39542),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_14_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_14_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_14_15_6  (
            .in0(N__44097),
            .in1(N__39114),
            .in2(_gnd_net_),
            .in3(N__42744),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(elapsed_time_ns_1_RNILK91B_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_14_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_14_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39108),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_14_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_14_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_0_LC_14_16_0  (
            .in0(N__39824),
            .in1(N__39086),
            .in2(N__39104),
            .in3(N__39105),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_0 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_14_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_14_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_1_LC_14_16_1  (
            .in0(N__39828),
            .in1(N__39071),
            .in2(_gnd_net_),
            .in3(N__39057),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_1 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_14_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_14_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_2_LC_14_16_2  (
            .in0(N__39825),
            .in1(N__39377),
            .in2(_gnd_net_),
            .in3(N__39363),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_2 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_14_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_14_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_3_LC_14_16_3  (
            .in0(N__39829),
            .in1(N__39359),
            .in2(_gnd_net_),
            .in3(N__39345),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_3 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_14_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_14_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_4_LC_14_16_4  (
            .in0(N__39826),
            .in1(N__39341),
            .in2(_gnd_net_),
            .in3(N__39327),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_4 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_14_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_14_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_5_LC_14_16_5  (
            .in0(N__39830),
            .in1(N__39323),
            .in2(_gnd_net_),
            .in3(N__39309),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_5 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_14_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_14_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_6_LC_14_16_6  (
            .in0(N__39827),
            .in1(N__39305),
            .in2(_gnd_net_),
            .in3(N__39291),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_6 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_14_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_14_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_7_LC_14_16_7  (
            .in0(N__39831),
            .in1(N__39287),
            .in2(_gnd_net_),
            .in3(N__39273),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_7 ),
            .clk(N__52423),
            .ce(N__39675),
            .sr(N__51958));
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_14_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_14_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_8_LC_14_17_0  (
            .in0(N__39811),
            .in1(N__39269),
            .in2(_gnd_net_),
            .in3(N__39255),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_8 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_14_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_14_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_9_LC_14_17_1  (
            .in0(N__39815),
            .in1(N__39251),
            .in2(_gnd_net_),
            .in3(N__39237),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_9 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_14_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_14_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_10_LC_14_17_2  (
            .in0(N__39808),
            .in1(N__39497),
            .in2(_gnd_net_),
            .in3(N__39483),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_10 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_14_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_14_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_11_LC_14_17_3  (
            .in0(N__39812),
            .in1(N__39479),
            .in2(_gnd_net_),
            .in3(N__39465),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_11 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_14_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_14_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_12_LC_14_17_4  (
            .in0(N__39809),
            .in1(N__39458),
            .in2(_gnd_net_),
            .in3(N__39444),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_12 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_14_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_14_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_13_LC_14_17_5  (
            .in0(N__39813),
            .in1(N__39440),
            .in2(_gnd_net_),
            .in3(N__39426),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_13 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_14_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_14_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_14_LC_14_17_6  (
            .in0(N__39810),
            .in1(N__39422),
            .in2(_gnd_net_),
            .in3(N__39408),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_14 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_14_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_14_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_15_LC_14_17_7  (
            .in0(N__39814),
            .in1(N__39404),
            .in2(_gnd_net_),
            .in3(N__39390),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_15 ),
            .clk(N__52418),
            .ce(N__39681),
            .sr(N__51964));
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_14_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_14_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_16_LC_14_18_0  (
            .in0(N__39800),
            .in1(N__41798),
            .in2(_gnd_net_),
            .in3(N__39387),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_16 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_14_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_14_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_17_LC_14_18_1  (
            .in0(N__39804),
            .in1(N__41825),
            .in2(_gnd_net_),
            .in3(N__39384),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_17 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_14_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_14_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_18_LC_14_18_2  (
            .in0(N__39801),
            .in1(N__41717),
            .in2(_gnd_net_),
            .in3(N__39381),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_18 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_14_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_14_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_19_LC_14_18_3  (
            .in0(N__39805),
            .in1(N__41744),
            .in2(_gnd_net_),
            .in3(N__39564),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_19 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_14_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_14_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_14_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_20_LC_14_18_4  (
            .in0(N__39802),
            .in1(N__41480),
            .in2(_gnd_net_),
            .in3(N__39561),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_20 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_14_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_14_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_21_LC_14_18_5  (
            .in0(N__39806),
            .in1(N__41501),
            .in2(_gnd_net_),
            .in3(N__39558),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_21 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_14_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_14_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_14_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_22_LC_14_18_6  (
            .in0(N__39803),
            .in1(N__41399),
            .in2(_gnd_net_),
            .in3(N__39555),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_22 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_14_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_14_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_23_LC_14_18_7  (
            .in0(N__39807),
            .in1(N__41426),
            .in2(_gnd_net_),
            .in3(N__39552),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_23 ),
            .clk(N__52412),
            .ce(N__39679),
            .sr(N__51967));
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_14_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_14_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_14_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_24_LC_14_19_0  (
            .in0(N__39816),
            .in1(N__41564),
            .in2(_gnd_net_),
            .in3(N__39549),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_24 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_14_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_14_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_14_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_25_LC_14_19_1  (
            .in0(N__39820),
            .in1(N__41605),
            .in2(_gnd_net_),
            .in3(N__39546),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_25 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_14_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_14_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_26_LC_14_19_2  (
            .in0(N__39817),
            .in1(N__39541),
            .in2(_gnd_net_),
            .in3(N__39525),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_26 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_14_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_14_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_27_LC_14_19_3  (
            .in0(N__39821),
            .in1(N__39515),
            .in2(_gnd_net_),
            .in3(N__39501),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_27 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_14_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_14_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_28_LC_14_19_4  (
            .in0(N__39818),
            .in1(N__39902),
            .in2(_gnd_net_),
            .in3(N__39888),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_28 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_14_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_14_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_29_LC_14_19_5  (
            .in0(N__39822),
            .in1(N__39875),
            .in2(_gnd_net_),
            .in3(N__39861),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_29 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_14_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_14_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_30_LC_14_19_6  (
            .in0(N__39819),
            .in1(N__39850),
            .in2(_gnd_net_),
            .in3(N__39834),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_30 ),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_14_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_14_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_31_LC_14_19_7  (
            .in0(N__39823),
            .in1(N__39697),
            .in2(_gnd_net_),
            .in3(N__39708),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52407),
            .ce(N__39680),
            .sr(N__51973));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_14_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_14_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__42281),
            .in2(N__39630),
            .in3(N__42197),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_14_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_14_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__39621),
            .in2(_gnd_net_),
            .in3(N__42104),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_14_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_14_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__42366),
            .in2(_gnd_net_),
            .in3(N__39582),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_14_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_14_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__43830),
            .in2(_gnd_net_),
            .in3(N__39567),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_14_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_14_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42447),
            .in3(N__40038),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_14_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_14_20_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42018),
            .in3(N__40023),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_14_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_14_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__42324),
            .in2(_gnd_net_),
            .in3(N__40008),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_14_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_14_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__42345),
            .in2(_gnd_net_),
            .in3(N__39993),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_14_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_14_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__39990),
            .in2(_gnd_net_),
            .in3(N__39960),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_14_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_14_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__42543),
            .in2(_gnd_net_),
            .in3(N__39942),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_14_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_14_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__41871),
            .in2(_gnd_net_),
            .in3(N__39927),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_14_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_14_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__41970),
            .in2(_gnd_net_),
            .in3(N__39912),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_14_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_14_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__42078),
            .in2(_gnd_net_),
            .in3(N__40188),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_14_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_14_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__42528),
            .in2(_gnd_net_),
            .in3(N__40173),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_14_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_14_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__43719),
            .in2(_gnd_net_),
            .in3(N__40158),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_14_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_14_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__42351),
            .in2(_gnd_net_),
            .in3(N__40143),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_14_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_14_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__41955),
            .in2(_gnd_net_),
            .in3(N__40122),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_14_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_14_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__42474),
            .in2(_gnd_net_),
            .in3(N__40104),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_14_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_14_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__43140),
            .in2(_gnd_net_),
            .in3(N__40089),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_14_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_14_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__42429),
            .in2(_gnd_net_),
            .in3(N__40068),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_14_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_14_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__42057),
            .in2(_gnd_net_),
            .in3(N__40053),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_14_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_14_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__42597),
            .in2(_gnd_net_),
            .in3(N__40317),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_14_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_14_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(N__42582),
            .in2(_gnd_net_),
            .in3(N__40302),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_14_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_14_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__42468),
            .in2(_gnd_net_),
            .in3(N__40287),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_14_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_14_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__42453),
            .in2(_gnd_net_),
            .in3(N__40266),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_14_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_14_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__41943),
            .in2(_gnd_net_),
            .in3(N__40248),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_14_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_14_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__42552),
            .in2(_gnd_net_),
            .in3(N__40233),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_14_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_14_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__42858),
            .in2(_gnd_net_),
            .in3(N__40218),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_14_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_14_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__42843),
            .in2(_gnd_net_),
            .in3(N__40203),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_14_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_14_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__42558),
            .in2(_gnd_net_),
            .in3(N__40482),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_14_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_14_23_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_14_23_6  (
            .in0(N__42294),
            .in1(N__40479),
            .in2(_gnd_net_),
            .in3(N__40473),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_24_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__40441),
            .in2(N__42230),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__40420),
            .in2(N__42182),
            .in3(N__40446),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__40442),
            .in2(N__40400),
            .in3(N__40428),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__40372),
            .in2(N__40425),
            .in3(N__40404),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(N__40348),
            .in2(N__40401),
            .in3(N__40380),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_24_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(N__40678),
            .in2(N__40377),
            .in3(N__40356),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_24_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_24_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__40654),
            .in2(N__40353),
            .in3(N__40332),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_24_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_24_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_24_7  (
            .in0(_gnd_net_),
            .in1(N__40633),
            .in2(N__40683),
            .in3(N__40662),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__52386),
            .ce(N__42147),
            .sr(N__52000));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_25_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_25_0  (
            .in0(_gnd_net_),
            .in1(N__40609),
            .in2(N__40659),
            .in3(N__40638),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_25_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_25_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(N__40635),
            .in2(N__40589),
            .in3(N__40617),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_25_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__40561),
            .in2(N__40614),
            .in3(N__40593),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_25_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_25_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(N__40537),
            .in2(N__40590),
            .in3(N__40569),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_25_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_25_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__40513),
            .in2(N__40566),
            .in3(N__40545),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_25_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_25_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__40864),
            .in2(N__40542),
            .in3(N__40521),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_25_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_25_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__40840),
            .in2(N__40518),
            .in3(N__40497),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_25_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_25_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__40816),
            .in2(N__40869),
            .in3(N__40848),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__52382),
            .ce(N__42157),
            .sr(N__52006));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__40795),
            .in2(N__40845),
            .in3(N__40824),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__40774),
            .in2(N__40821),
            .in3(N__40800),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__40796),
            .in2(N__40754),
            .in3(N__40782),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__40726),
            .in2(N__40779),
            .in3(N__40758),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__40702),
            .in2(N__40755),
            .in3(N__40734),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_26_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__41068),
            .in2(N__40731),
            .in3(N__40710),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_26_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_26_6  (
            .in0(_gnd_net_),
            .in1(N__41044),
            .in2(N__40707),
            .in3(N__40686),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_26_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_26_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(N__41023),
            .in2(N__41073),
            .in3(N__41052),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__52378),
            .ce(N__42159),
            .sr(N__52013));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_27_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_27_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_27_0  (
            .in0(_gnd_net_),
            .in1(N__40987),
            .in2(N__41049),
            .in3(N__41028),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__52375),
            .ce(N__42158),
            .sr(N__52022));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_27_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_27_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(N__41025),
            .in2(N__40955),
            .in3(N__41007),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__52375),
            .ce(N__42158),
            .sr(N__52022));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_27_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_27_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_27_2  (
            .in0(_gnd_net_),
            .in1(N__41003),
            .in2(N__40992),
            .in3(N__40971),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__52375),
            .ce(N__42158),
            .sr(N__52022));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_27_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_27_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_27_3  (
            .in0(_gnd_net_),
            .in1(N__40967),
            .in2(N__40956),
            .in3(N__40935),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__52375),
            .ce(N__42158),
            .sr(N__52022));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_27_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_27_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40932),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52375),
            .ce(N__42158),
            .sr(N__52022));
    defparam \phase_controller_inst1.S1_LC_14_29_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_14_29_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_14_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_14_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41229),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52371),
            .ce(),
            .sr(N__52035));
    defparam \current_shift_inst.timer_s1.running_LC_14_30_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_14_30_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_14_30_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_14_30_0  (
            .in0(N__41169),
            .in1(N__40921),
            .in2(_gnd_net_),
            .in3(N__40892),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52369),
            .ce(),
            .sr(N__52040));
    defparam \current_shift_inst.stop_timer_s1_LC_14_30_6 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_14_30_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_14_30_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_14_30_6  (
            .in0(N__41227),
            .in1(N__41243),
            .in2(N__41172),
            .in3(N__40891),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52369),
            .ce(),
            .sr(N__52040));
    defparam \current_shift_inst.start_timer_s1_LC_14_30_7 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_14_30_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_14_30_7 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_14_30_7  (
            .in0(N__41242),
            .in1(N__41170),
            .in2(_gnd_net_),
            .in3(N__41228),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52369),
            .ce(),
            .sr(N__52040));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_15_8_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_15_8_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_0_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__47643),
            .in2(_gnd_net_),
            .in3(N__47149),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52475),
            .ce(N__50147),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_15_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_3_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45722),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52475),
            .ce(N__50147),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_15_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_4_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45701),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52475),
            .ce(N__50147),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_15_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_15_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_1_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45764),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52475),
            .ce(N__50147),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_15_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_2_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45743),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52475),
            .ce(N__50147),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_15_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_15_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_6_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45935),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52475),
            .ce(N__50147),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45939),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52468),
            .ce(N__43456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_9_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__45900),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52468),
            .ce(N__43456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45834),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52468),
            .ce(N__43456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45768),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52468),
            .ce(N__43456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45852),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52468),
            .ce(N__43456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45747),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52468),
            .ce(N__43456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_10_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_10_0  (
            .in0(N__41331),
            .in1(N__41322),
            .in2(N__41301),
            .in3(N__41268),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_15_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_15_10_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_20_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__45992),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52463),
            .ce(N__50145),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_15_10_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_15_10_2  (
            .in0(N__41330),
            .in1(N__41321),
            .in2(N__41300),
            .in3(N__41267),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_15_10_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_15_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_21_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45975),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52463),
            .ce(N__50145),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_10_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_10_4  (
            .in0(N__41685),
            .in1(N__41664),
            .in2(N__41655),
            .in3(N__45789),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_15_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_22_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46940),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52463),
            .ce(N__50145),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_15_10_6 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_15_10_6  (
            .in0(N__41684),
            .in1(N__41663),
            .in2(N__41654),
            .in3(N__45788),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_15_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_15_11_0 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_15_11_0  (
            .in0(N__41616),
            .in1(N__43499),
            .in2(N__41582),
            .in3(N__43484),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_12_0 .LUT_INIT=16'b0000101010001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_15_12_0  (
            .in0(N__43560),
            .in1(N__41523),
            .in2(N__41513),
            .in3(N__41487),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_15_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_15_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_20_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45996),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52453),
            .ce(N__43468),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_15_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_15_12_2 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_15_12_2  (
            .in0(N__43559),
            .in1(N__41522),
            .in2(N__41514),
            .in3(N__41486),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_12_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_15_12_4  (
            .in0(N__41442),
            .in1(N__41433),
            .in2(N__41411),
            .in3(N__41847),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_15_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_22_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46944),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52453),
            .ce(N__43468),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_15_12_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_15_12_6  (
            .in0(N__41441),
            .in1(N__41432),
            .in2(N__41412),
            .in3(N__41846),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_15_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_23_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46923),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52453),
            .ce(N__43468),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_15_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_15_13_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_15_13_0  (
            .in0(N__43539),
            .in1(N__41832),
            .in2(N__41811),
            .in3(N__41775),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_15_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_15_13_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_15_13_2  (
            .in0(N__43538),
            .in1(N__41831),
            .in2(N__41810),
            .in3(N__41774),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_15_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_17_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49923),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52446),
            .ce(N__43470),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_15_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_15_13_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_15_13_4  (
            .in0(N__41760),
            .in1(N__41751),
            .in2(N__41730),
            .in3(N__43527),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_15_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_15_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_18_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49578),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52446),
            .ce(N__43470),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_15_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_15_13_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_15_13_6  (
            .in0(N__41759),
            .in1(N__41750),
            .in2(N__41729),
            .in3(N__43526),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_14_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_14_0  (
            .in0(N__50343),
            .in1(N__41691),
            .in2(_gnd_net_),
            .in3(N__50822),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(elapsed_time_ns_1_RNIK63T9_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_15_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_15_14_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41910),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_14_2  (
            .in0(N__41907),
            .in1(N__48090),
            .in2(_gnd_net_),
            .in3(N__50825),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_15_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_15_14_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41901),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_14_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_14_4  (
            .in0(N__41898),
            .in1(N__47916),
            .in2(_gnd_net_),
            .in3(N__50824),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_15_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_15_14_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41892),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_15_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_15_14_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_15_14_6  (
            .in0(N__41889),
            .in1(N__47868),
            .in2(_gnd_net_),
            .in3(N__50823),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(elapsed_time_ns_1_RNIL73T9_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_15_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_15_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41883),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_15_0  (
            .in0(N__41880),
            .in1(N__42807),
            .in2(_gnd_net_),
            .in3(N__44098),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_15_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_15_15_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41874),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_15_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_15_4  (
            .in0(N__41988),
            .in1(N__47937),
            .in2(_gnd_net_),
            .in3(N__50836),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(elapsed_time_ns_1_RNI68CN9_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_15_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_15_15_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41982),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_15_7  (
            .in0(N__50837),
            .in1(N__43659),
            .in2(_gnd_net_),
            .in3(N__48063),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_16_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_16_2  (
            .in0(N__41979),
            .in1(N__42768),
            .in2(_gnd_net_),
            .in3(N__44099),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(elapsed_time_ns_1_RNIV8OBB_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_15_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_15_16_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41973),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_15_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_15_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41930),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_15_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_15_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42044),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_17_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_17_1  (
            .in0(N__44071),
            .in1(N__41931),
            .in2(_gnd_net_),
            .in3(N__42672),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_17_2  (
            .in0(N__42702),
            .in1(N__41919),
            .in2(_gnd_net_),
            .in3(N__44069),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_15_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_15_17_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41913),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_15_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_15_17_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_15_17_4  (
            .in0(N__42872),
            .in1(N__42918),
            .in2(_gnd_net_),
            .in3(N__44073),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_15_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_15_17_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_15_17_5  (
            .in0(N__44070),
            .in1(N__42066),
            .in2(_gnd_net_),
            .in3(N__43110),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_15_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_15_17_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42060),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_15_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_15_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_15_17_7  (
            .in0(N__44072),
            .in1(N__42045),
            .in2(_gnd_net_),
            .in3(N__42957),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_15_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_15_18_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_15_18_1  (
            .in0(N__44264),
            .in1(N__42240),
            .in2(N__42006),
            .in3(N__42819),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_18_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_15_18_2  (
            .in0(N__42314),
            .in1(N__42681),
            .in2(N__42033),
            .in3(N__43047),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_15_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_15_18_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__42027),
            .in2(N__42030),
            .in3(N__42837),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(elapsed_time_ns_1_RNIIH91B_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_15_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_15_18_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42021),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_15_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_15_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_15_18_5  (
            .in0(N__42005),
            .in1(N__42333),
            .in2(_gnd_net_),
            .in3(N__44043),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(elapsed_time_ns_1_RNIJI91B_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_15_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_15_18_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42327),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_15_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_15_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_15_18_7  (
            .in0(N__42280),
            .in1(N__42315),
            .in2(_gnd_net_),
            .in3(N__44044),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_19_0  (
            .in0(N__42092),
            .in1(N__42113),
            .in2(N__43862),
            .in3(N__42206),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42234),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52413),
            .ce(N__42135),
            .sr(N__51968));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_19_2  (
            .in0(N__42198),
            .in1(N__42207),
            .in2(_gnd_net_),
            .in3(N__44092),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42186),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52413),
            .ce(N__42135),
            .sr(N__51968));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_19_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_19_4  (
            .in0(N__42105),
            .in1(N__42114),
            .in2(_gnd_net_),
            .in3(N__44093),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_19_5  (
            .in0(N__44094),
            .in1(N__42378),
            .in2(_gnd_net_),
            .in3(N__42093),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_15_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_15_20_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__44279),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_20_1  (
            .in0(N__44104),
            .in1(N__42438),
            .in2(_gnd_net_),
            .in3(N__43128),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_15_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_15_20_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42432),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_20_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_20_3  (
            .in0(N__42417),
            .in1(N__44444),
            .in2(_gnd_net_),
            .in3(N__44348),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_156_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_15_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_15_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42377),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_20_5  (
            .in0(N__44103),
            .in1(N__42360),
            .in2(_gnd_net_),
            .in3(N__42651),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_15_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_15_20_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42354),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_15_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_15_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44240),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_15_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_15_21_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_15_21_0  (
            .in0(N__42339),
            .in1(N__42786),
            .in2(_gnd_net_),
            .in3(N__44100),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_15_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_15_21_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42546),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_21_3  (
            .in0(N__44101),
            .in1(N__42723),
            .in2(_gnd_net_),
            .in3(N__42537),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_15_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_15_21_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42531),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_15_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_15_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_15_21_5  (
            .in0(N__42521),
            .in1(N__44552),
            .in2(N__44510),
            .in3(N__42504),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_15_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_15_21_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_15_21_6  (
            .in0(N__42483),
            .in1(N__42630),
            .in2(_gnd_net_),
            .in3(N__44102),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_15_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_15_21_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42477),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_15_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_15_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42575),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_15_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_15_22_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_15_22_1  (
            .in0(N__42462),
            .in1(N__44109),
            .in2(_gnd_net_),
            .in3(N__42939),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_15_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_15_22_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42456),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_15_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_15_22_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_15_22_3  (
            .in0(N__42606),
            .in1(N__43074),
            .in2(_gnd_net_),
            .in3(N__44107),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_15_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_15_22_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42600),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_15_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_15_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_15_22_5  (
            .in0(N__42591),
            .in1(N__43038),
            .in2(_gnd_net_),
            .in3(N__44108),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_15_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_15_22_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42585),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_15_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_15_22_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_15_22_7  (
            .in0(N__42576),
            .in1(N__43002),
            .in2(_gnd_net_),
            .in3(N__44110),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_15_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_15_23_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_15_23_0  (
            .in0(N__44112),
            .in1(N__42567),
            .in2(_gnd_net_),
            .in3(N__42981),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_15_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_15_23_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42561),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_15_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_15_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43968),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_15_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_15_23_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_15_23_3  (
            .in0(N__45011),
            .in1(N__45406),
            .in2(_gnd_net_),
            .in3(N__44949),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_15_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_15_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42876),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_15_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_15_23_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_15_23_5  (
            .in0(N__42852),
            .in1(N__43020),
            .in2(_gnd_net_),
            .in3(N__44111),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_15_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_15_23_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42846),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_15_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_15_23_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_15_23_7  (
            .in0(N__42830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44291),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_15_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_15_24_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_15_24_0  (
            .in0(N__42797),
            .in1(N__42779),
            .in2(N__42761),
            .in3(N__42734),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_15_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_15_24_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__42716),
            .in2(N__42705),
            .in3(N__42692),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_15_25_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_15_25_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_15_25_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_15_25_1  (
            .in0(N__42662),
            .in1(N__42641),
            .in2(N__43745),
            .in3(N__42623),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_15_25_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_15_25_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_15_25_2  (
            .in0(N__42612),
            .in1(N__43088),
            .in2(_gnd_net_),
            .in3(N__44106),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_15_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_15_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_15_25_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43143),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_15_26_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_15_26_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_15_26_0  (
            .in0(N__43121),
            .in1(N__43100),
            .in2(N__43089),
            .in3(N__43067),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_15_26_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_15_26_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_15_26_1  (
            .in0(N__43056),
            .in1(N__42963),
            .in2(N__43050),
            .in3(N__42897),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_15_26_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_15_26_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_15_26_3  (
            .in0(N__43031),
            .in1(N__43013),
            .in2(N__42998),
            .in3(N__42974),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_15_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_15_26_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_15_26_4  (
            .in0(N__44123),
            .in1(N__42950),
            .in2(N__42935),
            .in3(N__42908),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_15_27_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_15_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_15_27_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_15_27_6  (
            .in0(N__51149),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44711),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_28_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_15_28_0  (
            .in0(_gnd_net_),
            .in1(N__51300),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_28_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_15_28_1  (
            .in0(_gnd_net_),
            .in1(N__42891),
            .in2(_gnd_net_),
            .in3(N__42879),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_15_28_2  (
            .in0(_gnd_net_),
            .in1(N__43191),
            .in2(_gnd_net_),
            .in3(N__43176),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_15_28_3  (
            .in0(_gnd_net_),
            .in1(N__43173),
            .in2(_gnd_net_),
            .in3(N__43161),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_28_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_15_28_4  (
            .in0(_gnd_net_),
            .in1(N__44784),
            .in2(_gnd_net_),
            .in3(N__43158),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_28_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_28_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_15_28_5  (
            .in0(_gnd_net_),
            .in1(N__46829),
            .in2(N__45315),
            .in3(N__43155),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_28_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_28_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_15_28_6  (
            .in0(_gnd_net_),
            .in1(N__45261),
            .in2(N__46880),
            .in3(N__43152),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_28_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_28_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_15_28_7  (
            .in0(_gnd_net_),
            .in1(N__45213),
            .in2(N__46881),
            .in3(N__43149),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_29_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_29_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_15_29_0  (
            .in0(_gnd_net_),
            .in1(N__45174),
            .in2(_gnd_net_),
            .in3(N__43146),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_15_29_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_29_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_29_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_29_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_15_29_1  (
            .in0(_gnd_net_),
            .in1(N__45132),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_29_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_29_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_29_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_15_29_2  (
            .in0(_gnd_net_),
            .in1(N__45087),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_29_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_29_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_29_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_15_29_3  (
            .in0(_gnd_net_),
            .in1(N__45039),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_29_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_29_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_29_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_15_29_4  (
            .in0(_gnd_net_),
            .in1(N__45642),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_29_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_29_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_29_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_15_29_5  (
            .in0(_gnd_net_),
            .in1(N__45591),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_29_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_29_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_29_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_15_29_6  (
            .in0(_gnd_net_),
            .in1(N__45561),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_29_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_29_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_29_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_15_29_7  (
            .in0(_gnd_net_),
            .in1(N__45531),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_30_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_30_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_30_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_15_30_0  (
            .in0(_gnd_net_),
            .in1(N__45507),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_30_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_30_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_30_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_30_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_15_30_1  (
            .in0(_gnd_net_),
            .in1(N__45480),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_30_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_30_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_30_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_15_30_2  (
            .in0(_gnd_net_),
            .in1(N__45450),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_30_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_30_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_30_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_15_30_3  (
            .in0(_gnd_net_),
            .in1(N__45363),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_30_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_30_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_15_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43272),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_16_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_16_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_11_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45851),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52480),
            .ce(N__50146),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_16_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_16_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_14_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46038),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52480),
            .ce(N__50146),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_16_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_16_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_5_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45953),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52480),
            .ce(N__50146),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_16_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_16_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_7_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45914),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52480),
            .ce(N__50146),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_16_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_16_9_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_16_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_10_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45866),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52476),
            .ce(N__50131),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_16_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_16_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_15_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46022),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52476),
            .ce(N__50131),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_16_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_16_9_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_16_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_12_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45830),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52476),
            .ce(N__50131),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_16_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_16_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_9_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45881),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52476),
            .ce(N__50131),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_16_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_16_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_13_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46052),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52476),
            .ce(N__50131),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_16_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_16_9_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_16_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_8_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45896),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52476),
            .ce(N__50131),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_16_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_16_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_3_LC_16_10_0  (
            .in0(N__45723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_10_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46023),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_16_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_16_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_5_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45957),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_16_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_16_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_13_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46053),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_16_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_16_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_14_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46037),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_16_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_16_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_27_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50246),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_16_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_16_10_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_9_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__45882),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_16_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_16_10_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_16_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_10_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45867),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52469),
            .ce(N__43435),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_16_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_16_11_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_16_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_26_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50225),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_16_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_16_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_21_LC_16_11_1  (
            .in0(N__45974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_16_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_16_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_4_LC_16_11_2  (
            .in0(N__45702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_16_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_16_11_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_16_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__49589),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_16_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_16_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_19_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50015),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_16_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_16_11_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_16_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_7_LC_16_11_5  (
            .in0(N__45918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_16_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_16_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_24_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50204),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_16_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_25_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50183),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52464),
            .ce(N__43469),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_16_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_16_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_16_12_1  (
            .in0(N__43674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_12_2  (
            .in0(N__43611),
            .in1(N__47961),
            .in2(_gnd_net_),
            .in3(N__50847),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(elapsed_time_ns_1_RNI57CN9_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_16_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_16_12_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43605),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_12_6  (
            .in0(N__50715),
            .in1(N__43602),
            .in2(_gnd_net_),
            .in3(N__50846),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(elapsed_time_ns_1_RNIF13T9_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_16_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_16_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43596),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_13_0  (
            .in0(N__50325),
            .in1(N__43593),
            .in2(_gnd_net_),
            .in3(N__50850),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_16_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_16_13_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43587),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_16_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_16_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_16_13_2  (
            .in0(N__46095),
            .in1(N__50646),
            .in2(_gnd_net_),
            .in3(N__50848),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_13_3  (
            .in0(N__50849),
            .in1(N__46073),
            .in2(_gnd_net_),
            .in3(N__50601),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_13_4  (
            .in0(N__43584),
            .in1(N__48000),
            .in2(_gnd_net_),
            .in3(N__50852),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(elapsed_time_ns_1_RNI35CN9_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_13_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43647),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_16_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_16_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_16_13_6  (
            .in0(N__43644),
            .in1(N__47847),
            .in2(_gnd_net_),
            .in3(N__50851),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_16_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_16_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43638),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_16_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_16_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43703),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_14_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_14_1  (
            .in0(N__50697),
            .in1(N__43635),
            .in2(_gnd_net_),
            .in3(N__50815),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(elapsed_time_ns_1_RNIG23T9_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_16_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_16_14_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43629),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_14_3  (
            .in0(N__43626),
            .in1(N__48018),
            .in2(_gnd_net_),
            .in3(N__50817),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(elapsed_time_ns_1_RNI24CN9_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_16_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_16_14_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43620),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_14_5  (
            .in0(N__43617),
            .in1(N__48039),
            .in2(_gnd_net_),
            .in3(N__50816),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(elapsed_time_ns_1_RNI13CN9_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_16_14_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43707),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_14_7  (
            .in0(N__43704),
            .in1(N__48144),
            .in2(_gnd_net_),
            .in3(N__50818),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_16_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_16_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_16_15_0  (
            .in0(N__43695),
            .in1(N__47826),
            .in2(_gnd_net_),
            .in3(N__50833),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_16_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_16_15_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43689),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_16_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_16_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_16_15_2  (
            .in0(N__47979),
            .in1(N__43686),
            .in2(_gnd_net_),
            .in3(N__50834),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_16_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_16_15_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43680),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_16_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_16_15_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_16_15_4  (
            .in0(N__43785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_15_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_15_5  (
            .in0(N__43758),
            .in1(N__50907),
            .in2(N__43881),
            .in3(N__48326),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_16_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_16_15_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_16_15_6  (
            .in0(N__43673),
            .in1(_gnd_net_),
            .in2(N__43677),
            .in3(N__50370),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_16_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_16_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43658),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_16_0  (
            .in0(N__43770),
            .in1(N__48168),
            .in2(_gnd_net_),
            .in3(N__50845),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_16_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_16_16_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43764),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_16_5  (
            .in0(N__47822),
            .in1(N__47840),
            .in2(N__50057),
            .in3(N__47861),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_16_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__48032),
            .in2(N__43761),
            .in3(N__50426),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_16_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_16_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43800),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_17_0  (
            .in0(N__43752),
            .in1(N__43728),
            .in2(_gnd_net_),
            .in3(N__44074),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(elapsed_time_ns_1_RNI2COBB_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_16_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_16_17_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43722),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_17_4  (
            .in0(N__47975),
            .in1(N__47993),
            .in2(N__47957),
            .in3(N__48014),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_16_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43811),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_17_6  (
            .in0(N__47894),
            .in1(N__47909),
            .in2(N__48167),
            .in3(N__47930),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_16_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_16_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_16_17_7  (
            .in0(N__43890),
            .in1(N__43869),
            .in2(N__43884),
            .in3(N__43818),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_18_0  (
            .in0(N__50396),
            .in1(N__48104),
            .in2(N__48123),
            .in3(N__48080),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_18_1  (
            .in0(N__43863),
            .in1(N__43839),
            .in2(_gnd_net_),
            .in3(N__44042),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(elapsed_time_ns_1_RNIGF91B_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_16_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_16_18_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43833),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_18_3  (
            .in0(N__50891),
            .in1(N__48137),
            .in2(N__48059),
            .in3(N__50477),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_18_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_18_4  (
            .in0(N__43812),
            .in1(N__48105),
            .in2(_gnd_net_),
            .in3(N__50873),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_18_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__48122),
            .in2(N__50880),
            .in3(N__43799),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_18_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_18_6  (
            .in0(N__47895),
            .in1(N__43784),
            .in2(_gnd_net_),
            .in3(N__50869),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__44448),
            .in2(_gnd_net_),
            .in3(N__44349),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_155_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_19_1  (
            .in0(N__44280),
            .in1(N__44301),
            .in2(_gnd_net_),
            .in3(N__44095),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_19_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_19_3  (
            .in0(N__44241),
            .in1(N__44268),
            .in2(_gnd_net_),
            .in3(N__44096),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_16_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_16_20_1  (
            .in0(N__44229),
            .in1(N__44201),
            .in2(N__44181),
            .in3(N__44153),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_20_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_20_6  (
            .in0(N__43967),
            .in1(N__44133),
            .in2(_gnd_net_),
            .in3(N__44105),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_16_20_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_16_20_7  (
            .in0(N__44648),
            .in1(N__43952),
            .in2(N__44604),
            .in3(N__43931),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_16_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_16_21_0  (
            .in0(N__44565),
            .in1(N__43911),
            .in2(N__44538),
            .in3(N__44577),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_16_21_1  (
            .in0(N__43905),
            .in1(N__43899),
            .in2(N__43893),
            .in3(N__44355),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_16_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_16_21_2  (
            .in0(N__44603),
            .in1(N__44409),
            .in2(N__44388),
            .in3(N__44576),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_16_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_16_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__44564),
            .in2(_gnd_net_),
            .in3(N__44553),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_16_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_16_22_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__44528),
            .in2(_gnd_net_),
            .in3(N__44486),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_16_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_16_22_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_16_22_1  (
            .in0(N__44529),
            .in1(N__44514),
            .in2(N__44490),
            .in3(N__44475),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_2  (
            .in0(N__44634),
            .in1(N__44469),
            .in2(N__44463),
            .in3(N__44460),
            .lcout(\current_shift_inst.PI_CTRL.N_150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44437),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_16_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_16_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__44402),
            .in2(_gnd_net_),
            .in3(N__44387),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_16_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_16_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_16_22_6  (
            .in0(N__44687),
            .in1(N__44669),
            .in2(N__44358),
            .in3(N__44699),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_16_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_16_22_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_16_22_7  (
            .in0(N__44700),
            .in1(N__44688),
            .in2(N__44673),
            .in3(N__44655),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_16_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_16_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_16_23_0  (
            .in0(N__44757),
            .in1(N__48854),
            .in2(_gnd_net_),
            .in3(N__44628),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_1_LC_16_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_16_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_16_23_1  (
            .in0(N__44753),
            .in1(N__48827),
            .in2(_gnd_net_),
            .in3(N__44625),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_2_LC_16_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_16_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_16_23_2  (
            .in0(N__44758),
            .in1(N__49382),
            .in2(_gnd_net_),
            .in3(N__44622),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_3_LC_16_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_16_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_16_23_3  (
            .in0(N__44754),
            .in1(N__49355),
            .in2(_gnd_net_),
            .in3(N__44619),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_4_LC_16_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_16_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_16_23_4  (
            .in0(N__44759),
            .in1(N__49328),
            .in2(_gnd_net_),
            .in3(N__44616),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_5_LC_16_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_16_23_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_16_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_16_23_5  (
            .in0(N__44755),
            .in1(N__49301),
            .in2(_gnd_net_),
            .in3(N__44613),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_6_LC_16_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_16_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_16_23_6  (
            .in0(N__44760),
            .in1(N__49271),
            .in2(_gnd_net_),
            .in3(N__44610),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_7_LC_16_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_16_23_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_16_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_16_23_7  (
            .in0(N__44756),
            .in1(N__49247),
            .in2(_gnd_net_),
            .in3(N__44607),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__52399),
            .ce(),
            .sr(N__51978));
    defparam \pwm_generator_inst.counter_8_LC_16_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_16_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_16_24_0  (
            .in0(N__44752),
            .in1(N__49221),
            .in2(_gnd_net_),
            .in3(N__44778),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__52394),
            .ce(),
            .sr(N__51987));
    defparam \pwm_generator_inst.counter_9_LC_16_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_16_24_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_16_24_1  (
            .in0(N__49197),
            .in1(N__44751),
            .in2(_gnd_net_),
            .in3(N__44775),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52394),
            .ce(),
            .sr(N__51987));
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_16_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_16_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_16_25_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNITBL3_9_LC_16_25_1  (
            .in0(N__49219),
            .in1(N__49195),
            .in2(_gnd_net_),
            .in3(N__49302),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_16_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_16_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIRPD2_0_LC_16_25_5  (
            .in0(_gnd_net_),
            .in1(N__48855),
            .in2(_gnd_net_),
            .in3(N__48828),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_16_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_16_25_6 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_2_LC_16_25_6  (
            .in0(N__49329),
            .in1(N__49356),
            .in2(N__44772),
            .in3(N__49383),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_16_25_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_16_25_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_6_LC_16_25_7  (
            .in0(N__44769),
            .in1(N__49248),
            .in2(N__44763),
            .in3(N__49275),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_16_26_2  (
            .in0(N__51148),
            .in1(N__51369),
            .in2(N__44718),
            .in3(N__51129),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_16_26_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_16_26_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_16_26_3  (
            .in0(N__51426),
            .in1(N__51393),
            .in2(N__51379),
            .in3(N__51450),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_16_26_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_16_26_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_16_26_4  (
            .in0(N__51261),
            .in1(N__51234),
            .in2(N__44841),
            .in3(N__51367),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_16_26_5  (
            .in0(_gnd_net_),
            .in1(N__49640),
            .in2(_gnd_net_),
            .in3(N__51191),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_16_26_6  (
            .in0(_gnd_net_),
            .in1(N__51221),
            .in2(_gnd_net_),
            .in3(N__45026),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_16_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_16_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_16_26_7 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_16_26_7  (
            .in0(N__51368),
            .in1(N__51204),
            .in2(N__45030),
            .in3(N__45027),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_27_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_27_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_16_27_0  (
            .in0(N__49610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51496),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_16_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_16_27_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_16_27_1  (
            .in0(N__45012),
            .in1(N__45441),
            .in2(N__44979),
            .in3(N__44871),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_16_27_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_16_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_16_27_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_16_27_3  (
            .in0(_gnd_net_),
            .in1(N__44852),
            .in2(_gnd_net_),
            .in3(N__51080),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_16_27_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_16_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_16_27_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_16_27_4  (
            .in0(N__44853),
            .in1(N__51370),
            .in2(N__44844),
            .in3(N__51066),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_16_27_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_16_27_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_16_27_5  (
            .in0(N__51115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49664),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_27_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_27_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_16_27_7  (
            .in0(_gnd_net_),
            .in1(N__44834),
            .in2(_gnd_net_),
            .in3(N__51253),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_16_28_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_16_28_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_16_28_0  (
            .in0(_gnd_net_),
            .in1(N__44823),
            .in2(N__44802),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_16_28_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_28_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_16_28_1  (
            .in0(_gnd_net_),
            .in1(N__45357),
            .in2(N__45336),
            .in3(N__45306),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_28_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_16_28_2  (
            .in0(_gnd_net_),
            .in1(N__45303),
            .in2(N__45282),
            .in3(N__45255),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_28_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_16_28_3  (
            .in0(_gnd_net_),
            .in1(N__45252),
            .in2(N__45234),
            .in3(N__45207),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_28_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_16_28_4  (
            .in0(_gnd_net_),
            .in1(N__45204),
            .in2(N__45189),
            .in3(N__45168),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_28_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_16_28_5  (
            .in0(_gnd_net_),
            .in1(N__45165),
            .in2(N__45150),
            .in3(N__45126),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_28_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_16_28_6  (
            .in0(_gnd_net_),
            .in1(N__45123),
            .in2(N__45102),
            .in3(N__45081),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_28_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_28_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_16_28_7  (
            .in0(_gnd_net_),
            .in1(N__45078),
            .in2(N__45057),
            .in3(N__45033),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_29_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_29_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_16_29_0  (
            .in0(_gnd_net_),
            .in1(N__45681),
            .in2(N__45660),
            .in3(N__45636),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_16_29_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_29_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_29_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_16_29_1  (
            .in0(_gnd_net_),
            .in1(N__45633),
            .in2(N__45612),
            .in3(N__45585),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_29_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_29_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_16_29_2  (
            .in0(_gnd_net_),
            .in1(N__45582),
            .in2(N__45438),
            .in3(N__45555),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_29_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_29_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_16_29_3  (
            .in0(_gnd_net_),
            .in1(N__45426),
            .in2(N__45552),
            .in3(N__45525),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_29_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_29_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_16_29_4  (
            .in0(_gnd_net_),
            .in1(N__45522),
            .in2(N__45439),
            .in3(N__45501),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_29_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_29_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_16_29_5  (
            .in0(_gnd_net_),
            .in1(N__45430),
            .in2(N__45498),
            .in3(N__45474),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_29_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_29_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_16_29_6  (
            .in0(_gnd_net_),
            .in1(N__45471),
            .in2(N__45440),
            .in3(N__45444),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_29_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_29_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_16_29_7  (
            .in0(_gnd_net_),
            .in1(N__45434),
            .in2(N__45378),
            .in3(N__45816),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_30_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_30_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_30_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_16_30_0  (
            .in0(N__45813),
            .in1(N__45807),
            .in2(_gnd_net_),
            .in3(N__45798),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_16_30_2.C_ON=1'b0;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_16_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_16_30_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_red_c_g_THRU_LUT4_0_LC_16_30_2 (
            .in0(N__52086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_red_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_17_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_17_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_23_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46922),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52489),
            .ce(N__50156),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_17_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_17_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__45774),
            .in2(N__47153),
            .in3(N__47635),
            .lcout(\phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_17_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_17_8_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_17_8_1  (
            .in0(N__47103),
            .in1(N__47102),
            .in2(N__46757),
            .in3(N__45750),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_1),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_17_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_17_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_17_8_2  (
            .in0(N__47082),
            .in1(N__47081),
            .in2(N__46761),
            .in3(N__45726),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_2),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_17_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_17_8_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_17_8_3  (
            .in0(N__47058),
            .in1(N__47057),
            .in2(N__46758),
            .in3(N__45705),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_3),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_17_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_17_8_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_17_8_4  (
            .in0(N__47034),
            .in1(N__47033),
            .in2(N__46762),
            .in3(N__45684),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_4),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_17_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_17_8_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_17_8_5  (
            .in0(N__47001),
            .in1(N__47000),
            .in2(N__46759),
            .in3(N__45942),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_5),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_17_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_17_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_17_8_6  (
            .in0(N__46968),
            .in1(N__46967),
            .in2(N__46763),
            .in3(N__45921),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_6),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_17_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_17_8_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_17_8_7  (
            .in0(N__47367),
            .in1(N__47363),
            .in2(N__46760),
            .in3(N__45903),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_7),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_17_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_17_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_17_9_0  (
            .in0(N__47334),
            .in1(N__47333),
            .in2(N__46852),
            .in3(N__45885),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_8),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_17_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_17_9_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_17_9_1  (
            .in0(N__47313),
            .in1(N__47312),
            .in2(N__46771),
            .in3(N__45870),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_9),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_17_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_17_9_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_17_9_2  (
            .in0(N__47292),
            .in1(N__47291),
            .in2(N__46853),
            .in3(N__45855),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_10),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_17_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_17_9_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_17_9_3  (
            .in0(N__47262),
            .in1(N__47261),
            .in2(N__46768),
            .in3(N__45837),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_11),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_17_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_17_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_17_9_4  (
            .in0(N__47235),
            .in1(N__47234),
            .in2(N__46850),
            .in3(N__45819),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_12),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_17_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_17_9_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_17_9_5  (
            .in0(N__47211),
            .in1(N__47210),
            .in2(N__46769),
            .in3(N__46041),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_13),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_17_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_17_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_17_9_6  (
            .in0(N__47181),
            .in1(N__47180),
            .in2(N__46851),
            .in3(N__46026),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_14),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_17_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_17_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_17_9_7  (
            .in0(N__47574),
            .in1(N__47573),
            .in2(N__46770),
            .in3(N__46011),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_15),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_17_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_17_10_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_17_10_0  (
            .in0(N__47541),
            .in1(N__47540),
            .in2(N__46882),
            .in3(N__46008),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_16),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_17_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_17_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_17_10_1  (
            .in0(N__47511),
            .in1(N__47510),
            .in2(N__46764),
            .in3(N__46005),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_17),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_17_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_17_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_17_10_2  (
            .in0(N__47484),
            .in1(N__47483),
            .in2(N__46883),
            .in3(N__46002),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_18),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_17_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_17_10_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_17_10_3  (
            .in0(N__47457),
            .in1(N__47456),
            .in2(N__46765),
            .in3(N__45999),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_19),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_17_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_17_10_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_17_10_4  (
            .in0(N__47436),
            .in1(N__47435),
            .in2(N__46884),
            .in3(N__45978),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_20),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_17_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_17_10_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_17_10_5  (
            .in0(N__47412),
            .in1(N__47411),
            .in2(N__46766),
            .in3(N__45960),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_21),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_17_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_17_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_17_10_6  (
            .in0(N__47388),
            .in1(N__47387),
            .in2(N__46885),
            .in3(N__46926),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_22),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_17_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_17_10_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_17_10_7  (
            .in0(N__47796),
            .in1(N__47795),
            .in2(N__46767),
            .in3(N__46899),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_23),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_17_11_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_17_11_0  (
            .in0(N__47775),
            .in1(N__47774),
            .in2(N__46886),
            .in3(N__46896),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_24),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_17_11_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_17_11_1  (
            .in0(N__47745),
            .in1(N__47744),
            .in2(N__46848),
            .in3(N__46893),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_25),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_17_11_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_17_11_2  (
            .in0(N__47727),
            .in1(N__47726),
            .in2(N__46887),
            .in3(N__46890),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_26),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_17_11_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_17_11_3  (
            .in0(N__47700),
            .in1(N__47699),
            .in2(N__46849),
            .in3(N__46101),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_27),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_17_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_17_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46098),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_17_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__47625),
            .in2(N__46083),
            .in3(N__46094),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_17_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__46059),
            .in2(_gnd_net_),
            .in3(N__46074),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_17_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__47163),
            .in2(_gnd_net_),
            .in3(N__47115),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_17_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_17_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__47112),
            .in2(_gnd_net_),
            .in3(N__47085),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_17_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_17_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__50025),
            .in2(_gnd_net_),
            .in3(N__47067),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_17_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_17_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__47064),
            .in2(_gnd_net_),
            .in3(N__47043),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_17_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_17_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__47040),
            .in2(_gnd_net_),
            .in3(N__47016),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_17_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_17_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__47013),
            .in2(_gnd_net_),
            .in3(N__46983),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_17_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_17_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__46980),
            .in2(_gnd_net_),
            .in3(N__46953),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_17_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_17_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__46950),
            .in2(_gnd_net_),
            .in3(N__47346),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_17_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_17_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__47343),
            .in2(_gnd_net_),
            .in3(N__47316),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_17_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_17_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__50031),
            .in2(_gnd_net_),
            .in3(N__47295),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_17_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_17_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__50436),
            .in2(_gnd_net_),
            .in3(N__47271),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_17_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_17_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__47268),
            .in2(_gnd_net_),
            .in3(N__47244),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_17_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_17_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__47241),
            .in2(_gnd_net_),
            .in3(N__47220),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_17_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_17_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__47217),
            .in2(_gnd_net_),
            .in3(N__47190),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_17_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_17_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__47187),
            .in2(_gnd_net_),
            .in3(N__47166),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_17_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_17_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__47583),
            .in2(_gnd_net_),
            .in3(N__47556),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_17_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_17_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__47553),
            .in2(_gnd_net_),
            .in3(N__47523),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_17_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_17_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__47520),
            .in2(_gnd_net_),
            .in3(N__47493),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_17_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_17_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__47490),
            .in2(_gnd_net_),
            .in3(N__47469),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_17_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_17_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__47466),
            .in2(_gnd_net_),
            .in3(N__47439),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_17_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_17_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__50457),
            .in2(_gnd_net_),
            .in3(N__47421),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_17_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_17_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__47418),
            .in2(_gnd_net_),
            .in3(N__47397),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_17_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_17_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__47394),
            .in2(_gnd_net_),
            .in3(N__47370),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_17_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_17_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__47805),
            .in2(_gnd_net_),
            .in3(N__47778),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_17_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_17_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__50376),
            .in2(_gnd_net_),
            .in3(N__47760),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_17_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_17_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__47757),
            .in2(_gnd_net_),
            .in3(N__47730),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_17_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_17_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__50721),
            .in2(_gnd_net_),
            .in3(N__47709),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_17_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_17_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__47706),
            .in2(_gnd_net_),
            .in3(N__47685),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_17_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_17_15_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_17_15_6  (
            .in0(N__47682),
            .in1(N__47617),
            .in2(_gnd_net_),
            .in3(N__47670),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_17_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_17_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_17_15_7  (
            .in0(N__47618),
            .in1(N__48327),
            .in2(_gnd_net_),
            .in3(N__50835),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_16_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__48299),
            .in2(N__50673),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__48278),
            .in2(N__50628),
            .in3(N__47586),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__48300),
            .in2(N__48258),
            .in3(N__47880),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__48279),
            .in2(N__48231),
            .in3(N__47877),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__48257),
            .in2(N__48197),
            .in3(N__47874),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__48230),
            .in2(N__48578),
            .in3(N__47871),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__48542),
            .in2(N__48198),
            .in3(N__47850),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__48512),
            .in2(N__48579),
            .in3(N__47829),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__52440),
            .ce(N__50582),
            .sr(N__51946));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__48485),
            .in2(N__48549),
            .in3(N__47811),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__48461),
            .in2(N__48516),
            .in3(N__47808),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__48486),
            .in2(N__48437),
            .in3(N__48042),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__48462),
            .in2(N__48407),
            .in3(N__48021),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__48377),
            .in2(N__48438),
            .in3(N__48003),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__48353),
            .in2(N__48408),
            .in3(N__47982),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__48378),
            .in2(N__48797),
            .in3(N__47964),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__48354),
            .in2(N__48765),
            .in3(N__47940),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__52435),
            .ce(N__50574),
            .sr(N__51952));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__48728),
            .in2(N__48798),
            .in3(N__47919),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__48764),
            .in2(N__48701),
            .in3(N__47898),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__48674),
            .in2(N__48732),
            .in3(N__47883),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__48650),
            .in2(N__48702),
            .in3(N__48150),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__48675),
            .in2(N__48626),
            .in3(N__48147),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__48599),
            .in2(N__48654),
            .in3(N__48126),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__49166),
            .in2(N__48627),
            .in3(N__48108),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__48600),
            .in2(N__49136),
            .in3(N__48096),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__52430),
            .ce(N__50573),
            .sr(N__51955));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__49103),
            .in2(N__49173),
            .in3(N__48093),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__52424),
            .ce(N__50575),
            .sr(N__51959));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__49082),
            .in2(N__49140),
            .in3(N__48069),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__52424),
            .ce(N__50575),
            .sr(N__51959));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__49104),
            .in2(N__49062),
            .in3(N__48066),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__52424),
            .ce(N__50575),
            .sr(N__51959));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__49083),
            .in2(N__48921),
            .in3(N__48333),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__52424),
            .ce(N__50575),
            .sr(N__51959));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48330),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52424),
            .ce(N__50575),
            .sr(N__51959));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_20_0  (
            .in0(N__49034),
            .in1(N__50662),
            .in2(_gnd_net_),
            .in3(N__48306),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_20_1  (
            .in0(N__49030),
            .in1(N__50617),
            .in2(_gnd_net_),
            .in3(N__48303),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_20_2  (
            .in0(N__49035),
            .in1(N__48298),
            .in2(_gnd_net_),
            .in3(N__48282),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_20_3  (
            .in0(N__49031),
            .in1(N__48277),
            .in2(_gnd_net_),
            .in3(N__48261),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_20_4  (
            .in0(N__49036),
            .in1(N__48253),
            .in2(_gnd_net_),
            .in3(N__48234),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_20_5  (
            .in0(N__49032),
            .in1(N__48220),
            .in2(_gnd_net_),
            .in3(N__48201),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_20_6  (
            .in0(N__49037),
            .in1(N__48185),
            .in2(_gnd_net_),
            .in3(N__48171),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_20_7  (
            .in0(N__49033),
            .in1(N__48566),
            .in2(_gnd_net_),
            .in3(N__48552),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__52419),
            .ce(N__48888),
            .sr(N__51965));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_21_0  (
            .in0(N__49019),
            .in1(N__48541),
            .in2(_gnd_net_),
            .in3(N__48519),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_21_1  (
            .in0(N__49041),
            .in1(N__48505),
            .in2(_gnd_net_),
            .in3(N__48489),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_21_2  (
            .in0(N__49016),
            .in1(N__48479),
            .in2(_gnd_net_),
            .in3(N__48465),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_21_3  (
            .in0(N__49038),
            .in1(N__48455),
            .in2(_gnd_net_),
            .in3(N__48441),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_21_4  (
            .in0(N__49017),
            .in1(N__48425),
            .in2(_gnd_net_),
            .in3(N__48411),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_21_5  (
            .in0(N__49039),
            .in1(N__48395),
            .in2(_gnd_net_),
            .in3(N__48381),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_21_6  (
            .in0(N__49018),
            .in1(N__48371),
            .in2(_gnd_net_),
            .in3(N__48357),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_21_7  (
            .in0(N__49040),
            .in1(N__48347),
            .in2(_gnd_net_),
            .in3(N__48801),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__52414),
            .ce(N__48898),
            .sr(N__51969));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_22_0  (
            .in0(N__49012),
            .in1(N__48784),
            .in2(_gnd_net_),
            .in3(N__48768),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_22_1  (
            .in0(N__49026),
            .in1(N__48754),
            .in2(_gnd_net_),
            .in3(N__48735),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_22_2  (
            .in0(N__49013),
            .in1(N__48721),
            .in2(_gnd_net_),
            .in3(N__48705),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_22_3  (
            .in0(N__49027),
            .in1(N__48694),
            .in2(_gnd_net_),
            .in3(N__48678),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_22_4  (
            .in0(N__49014),
            .in1(N__48673),
            .in2(_gnd_net_),
            .in3(N__48657),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_22_5  (
            .in0(N__49028),
            .in1(N__48649),
            .in2(_gnd_net_),
            .in3(N__48630),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_22_6  (
            .in0(N__49015),
            .in1(N__48619),
            .in2(_gnd_net_),
            .in3(N__48603),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_22_7  (
            .in0(N__49029),
            .in1(N__48598),
            .in2(_gnd_net_),
            .in3(N__48582),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__52408),
            .ce(N__48903),
            .sr(N__51974));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_23_0  (
            .in0(N__49020),
            .in1(N__49165),
            .in2(_gnd_net_),
            .in3(N__49143),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__52403),
            .ce(N__48902),
            .sr(N__51975));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_23_1  (
            .in0(N__49024),
            .in1(N__49129),
            .in2(_gnd_net_),
            .in3(N__49107),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__52403),
            .ce(N__48902),
            .sr(N__51975));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_23_2  (
            .in0(N__49021),
            .in1(N__49102),
            .in2(_gnd_net_),
            .in3(N__49086),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__52403),
            .ce(N__48902),
            .sr(N__51975));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_23_3  (
            .in0(N__49025),
            .in1(N__49081),
            .in2(_gnd_net_),
            .in3(N__49065),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__52403),
            .ce(N__48902),
            .sr(N__51975));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_23_4  (
            .in0(N__49022),
            .in1(N__49058),
            .in2(_gnd_net_),
            .in3(N__49044),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__52403),
            .ce(N__48902),
            .sr(N__51975));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_23_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_23_5  (
            .in0(N__48917),
            .in1(N__49023),
            .in2(_gnd_net_),
            .in3(N__48924),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52403),
            .ce(N__48902),
            .sr(N__51975));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_17_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_17_24_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_17_24_0  (
            .in0(N__48853),
            .in1(N__48834),
            .in2(N__49524),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_17_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_17_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__48807),
            .in2(N__49509),
            .in3(N__48826),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_17_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_17_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__49362),
            .in2(N__49482),
            .in3(N__49378),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_17_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_17_24_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_17_24_3  (
            .in0(N__49351),
            .in1(N__49335),
            .in2(N__49458),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_17_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_17_24_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_17_24_4  (
            .in0(N__49324),
            .in1(N__49308),
            .in2(N__49440),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_17_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_17_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_17_24_5  (
            .in0(_gnd_net_),
            .in1(N__49281),
            .in2(N__49419),
            .in3(N__49297),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_17_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_17_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(N__49254),
            .in2(N__49401),
            .in3(N__49270),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_17_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_17_24_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_17_24_7  (
            .in0(N__49243),
            .in1(N__49227),
            .in2(N__49731),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_17_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_17_25_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_17_25_0  (
            .in0(N__49220),
            .in1(N__49203),
            .in2(N__49713),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_17_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_17_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_17_25_1  (
            .in0(_gnd_net_),
            .in1(N__49179),
            .in2(N__49683),
            .in3(N__49196),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_17_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_17_25_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_17_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_17_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49557),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52395),
            .ce(),
            .sr(N__51988));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_17_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_17_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__49530),
            .in2(N__51381),
            .in3(N__51380),
            .lcout(\pwm_generator_inst.un14_counter_0 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_0_c_RNI2C682_LC_17_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_0_c_RNI2C682_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_0_c_RNI2C682_LC_17_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_0_c_RNI2C682_LC_17_26_1  (
            .in0(_gnd_net_),
            .in1(N__51273),
            .in2(_gnd_net_),
            .in3(N__49494),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_1_c_RNI93892_LC_17_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_1_c_RNI93892_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_1_c_RNI93892_LC_17_26_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_1_c_RNI93892_LC_17_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49491),
            .in3(N__49467),
            .lcout(\pwm_generator_inst.un14_counter_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_2_c_RNIC9B92_LC_17_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_2_c_RNIC9B92_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_2_c_RNIC9B92_LC_17_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_2_c_RNIC9B92_LC_17_26_3  (
            .in0(_gnd_net_),
            .in1(N__49464),
            .in2(_gnd_net_),
            .in3(N__49443),
            .lcout(\pwm_generator_inst.un14_counter_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_3_c_RNIFFE92_LC_17_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_3_c_RNIFFE92_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_3_c_RNIFFE92_LC_17_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_3_c_RNIFFE92_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__49623),
            .in2(_gnd_net_),
            .in3(N__49428),
            .lcout(\pwm_generator_inst.un14_counter_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_4_c_RNI0V9N2_LC_17_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_4_c_RNI0V9N2_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_4_c_RNI0V9N2_LC_17_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_4_c_RNI0V9N2_LC_17_26_5  (
            .in0(_gnd_net_),
            .in1(N__49425),
            .in2(_gnd_net_),
            .in3(N__49404),
            .lcout(\pwm_generator_inst.un14_counter_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_5_c_RNIVCMU2_LC_17_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_5_c_RNIVCMU2_LC_17_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_5_c_RNIVCMU2_LC_17_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_5_c_RNIVCMU2_LC_17_26_6  (
            .in0(_gnd_net_),
            .in1(N__49653),
            .in2(_gnd_net_),
            .in3(N__49386),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_6_c_RNI3LQU2_LC_17_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_6_c_RNI3LQU2_LC_17_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_6_c_RNI3LQU2_LC_17_26_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_6_c_RNI3LQU2_LC_17_26_7  (
            .in0(_gnd_net_),
            .in1(N__49737),
            .in2(_gnd_net_),
            .in3(N__49716),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_0_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_0_cry_7_c_RNI7TUU2_LC_17_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_0_cry_7_c_RNI7TUU2_LC_17_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_0_cry_7_c_RNI7TUU2_LC_17_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_0_cry_7_c_RNI7TUU2_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(N__49599),
            .in2(_gnd_net_),
            .in3(N__49701),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(bfn_17_27_0_),
            .carryout(\pwm_generator_inst.un19_threshold_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIB53V2_LC_17_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIB53V2_LC_17_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIB53V2_LC_17_27_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIB53V2_LC_17_27_1  (
            .in0(N__51459),
            .in1(N__49698),
            .in2(N__51378),
            .in3(N__49686),
            .lcout(\pwm_generator_inst.un14_counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_17_27_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_17_27_4 .LUT_INIT=16'b1011011110000100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_17_27_4  (
            .in0(N__51093),
            .in1(N__51359),
            .in2(N__51117),
            .in3(N__49671),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_17_27_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_17_27_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_17_27_6  (
            .in0(N__51171),
            .in1(N__51190),
            .in2(N__49647),
            .in3(N__51358),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_17_27_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_17_27_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_17_27_7 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_17_27_7  (
            .in0(N__51360),
            .in1(N__49617),
            .in2(N__51498),
            .in3(N__51474),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_18_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_18_8_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_18_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_16_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49593),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52490),
            .ce(N__50141),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_18_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_18_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_18_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49577),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52490),
            .ce(N__50141),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_18_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_18_8_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_18_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_19_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50019),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52490),
            .ce(N__50141),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_18_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_18_9_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_18_9_0  (
            .in0(N__49992),
            .in1(N__49982),
            .in2(N__49964),
            .in3(N__49905),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_18_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_18_9_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_18_9_2  (
            .in0(N__49991),
            .in1(N__49983),
            .in2(N__49965),
            .in3(N__49904),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_18_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_18_9_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_18_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_17_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49916),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52484),
            .ce(N__50157),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_18_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_18_9_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_18_9_4  (
            .in0(N__49881),
            .in1(N__49872),
            .in2(N__49850),
            .in3(N__49827),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_18_9_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_18_9_6  (
            .in0(N__49880),
            .in1(N__49871),
            .in2(N__49851),
            .in3(N__49826),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_18_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_18_10_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_18_10_0  (
            .in0(N__50193),
            .in1(N__49791),
            .in2(N__50172),
            .in3(N__49773),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_18_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_18_10_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_18_10_2  (
            .in0(N__50192),
            .in1(N__49790),
            .in2(N__50171),
            .in3(N__49772),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_18_10_4 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_18_10_4  (
            .in0(N__50214),
            .in1(N__50307),
            .in2(N__50288),
            .in3(N__50235),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_18_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_18_10_6 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_18_10_6  (
            .in0(N__50213),
            .in1(N__50306),
            .in2(N__50289),
            .in3(N__50234),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_18_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_18_10_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_18_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_27_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50247),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52481),
            .ce(N__50140),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_18_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_18_11_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_18_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_26_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50226),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52477),
            .ce(N__50148),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_18_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_18_11_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_18_11_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_24_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__50205),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52477),
            .ce(N__50148),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_18_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_18_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_25_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50184),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52477),
            .ce(N__50148),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_18_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_18_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_18_12_0  (
            .in0(N__50040),
            .in1(N__50061),
            .in2(_gnd_net_),
            .in3(N__50875),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_18_12_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50034),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_18_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_18_12_3  (
            .in0(N__50447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_18_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_18_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_18_12_4  (
            .in0(N__50466),
            .in1(N__50484),
            .in2(_gnd_net_),
            .in3(N__50876),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(elapsed_time_ns_1_RNI14DN9_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_18_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_18_12_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50460),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_18_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_18_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_18_13_4  (
            .in0(N__50358),
            .in1(N__50448),
            .in2(_gnd_net_),
            .in3(N__50874),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_18_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_18_13_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__50414),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_14_0  (
            .in0(N__50877),
            .in1(N__50415),
            .in2(_gnd_net_),
            .in3(N__50430),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_14_5  (
            .in0(N__50385),
            .in1(N__50403),
            .in2(_gnd_net_),
            .in3(N__50878),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(elapsed_time_ns_1_RNI58DN9_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_14_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50379),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_18_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_18_15_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__50369),
            .in2(_gnd_net_),
            .in3(N__50354),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_18_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_18_15_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_18_15_1  (
            .in0(N__50336),
            .in1(N__50321),
            .in2(N__50310),
            .in3(N__50679),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_18_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_18_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_18_15_2  (
            .in0(N__50730),
            .in1(N__50898),
            .in2(_gnd_net_),
            .in3(N__50879),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_18_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_18_15_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50724),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_18_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_18_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_18_15_4  (
            .in0(N__50708),
            .in1(N__50594),
            .in2(N__50696),
            .in3(N__50639),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50672),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52447),
            .ce(N__50583),
            .sr(N__51944));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50627),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52447),
            .ce(N__50583),
            .sr(N__51944));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_20_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_20_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_20_25_0  (
            .in0(_gnd_net_),
            .in1(N__50526),
            .in2(_gnd_net_),
            .in3(N__50541),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_20_25_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_20_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_20_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_20_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_20_25_1  (
            .in0(_gnd_net_),
            .in1(N__50508),
            .in2(_gnd_net_),
            .in3(N__50520),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_20_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_20_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_20_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_20_25_2  (
            .in0(_gnd_net_),
            .in1(N__50490),
            .in2(_gnd_net_),
            .in3(N__50502),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_20_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_20_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_20_25_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_20_25_3  (
            .in0(_gnd_net_),
            .in1(N__51036),
            .in2(_gnd_net_),
            .in3(N__51051),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_20_25_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_20_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_20_25_4  (
            .in0(_gnd_net_),
            .in1(N__51015),
            .in2(_gnd_net_),
            .in3(N__51030),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_20_25_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_20_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_20_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_20_25_5  (
            .in0(_gnd_net_),
            .in1(N__50994),
            .in2(_gnd_net_),
            .in3(N__51009),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_20_25_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_20_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_20_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_20_25_6  (
            .in0(_gnd_net_),
            .in1(N__50973),
            .in2(_gnd_net_),
            .in3(N__50988),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_20_25_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_20_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_20_25_7  (
            .in0(_gnd_net_),
            .in1(N__50952),
            .in2(_gnd_net_),
            .in3(N__50967),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_20_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_20_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_20_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_20_26_0  (
            .in0(_gnd_net_),
            .in1(N__50931),
            .in2(_gnd_net_),
            .in3(N__50946),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_20_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_20_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_20_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_20_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_20_26_1  (
            .in0(_gnd_net_),
            .in1(N__50913),
            .in2(_gnd_net_),
            .in3(N__50925),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_20_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_20_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_20_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_20_26_2  (
            .in0(_gnd_net_),
            .in1(N__51421),
            .in2(_gnd_net_),
            .in3(N__51384),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_20_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_20_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_20_26_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_20_26_3  (
            .in0(N__51374),
            .in1(N__51299),
            .in2(_gnd_net_),
            .in3(N__51264),
            .lcout(\pwm_generator_inst.un19_threshold_0_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_20_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_20_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_20_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_20_26_4  (
            .in0(_gnd_net_),
            .in1(N__51260),
            .in2(_gnd_net_),
            .in3(N__51225),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_20_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_20_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_20_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_20_26_5  (
            .in0(_gnd_net_),
            .in1(N__51222),
            .in2(_gnd_net_),
            .in3(N__51195),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_20_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_20_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_20_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_20_26_6  (
            .in0(_gnd_net_),
            .in1(N__51192),
            .in2(_gnd_net_),
            .in3(N__51159),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_20_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_20_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_20_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_20_26_7  (
            .in0(_gnd_net_),
            .in1(N__51156),
            .in2(_gnd_net_),
            .in3(N__51120),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_20_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_20_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_20_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_20_27_0  (
            .in0(_gnd_net_),
            .in1(N__51116),
            .in2(_gnd_net_),
            .in3(N__51084),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_20_27_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_20_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_20_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_20_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_20_27_1  (
            .in0(_gnd_net_),
            .in1(N__51081),
            .in2(_gnd_net_),
            .in3(N__51054),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_20_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_20_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_20_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_20_27_2  (
            .in0(_gnd_net_),
            .in1(N__51497),
            .in2(_gnd_net_),
            .in3(N__51465),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_20_27_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_20_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_20_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_20_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51462),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_21_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_21_22_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_21_22_6  (
            .in0(N__52726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52825),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_21_26_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_21_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_21_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_21_26_2  (
            .in0(N__51425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51449),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_21_2  (
            .in0(_gnd_net_),
            .in1(N__52774),
            .in2(_gnd_net_),
            .in3(N__52727),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_22_1  (
            .in0(N__52862),
            .in1(N__51405),
            .in2(N__52826),
            .in3(N__52532),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_22_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_22_22_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_22_22_2  (
            .in0(N__52531),
            .in1(N__52861),
            .in2(N__52781),
            .in3(N__51399),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_21_7  (
            .in0(_gnd_net_),
            .in1(N__52929),
            .in2(_gnd_net_),
            .in3(N__51562),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_22_1 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_22_1  (
            .in0(N__52625),
            .in1(N__51676),
            .in2(N__52939),
            .in3(N__52561),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_22_2 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_22_2  (
            .in0(N__51693),
            .in1(N__52626),
            .in2(N__52895),
            .in3(N__52672),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_22_3 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_22_3  (
            .in0(N__51563),
            .in1(N__51684),
            .in2(N__51687),
            .in3(N__51527),
            .lcout(\current_shift_inst.PI_CTRL.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_22_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_22_6  (
            .in0(N__51677),
            .in1(N__52560),
            .in2(_gnd_net_),
            .in3(N__52624),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_7 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_22_7  (
            .in0(N__52627),
            .in1(N__51678),
            .in2(N__52940),
            .in3(N__52562),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51666),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52454),
            .ce(),
            .sr(N__51979));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_24_22_1  (
            .in0(N__51606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51651),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52448),
            .ce(),
            .sr(N__51990));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_24_22_2  (
            .in0(N__51621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51604),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52448),
            .ce(),
            .sr(N__51990));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_24_22_5  (
            .in0(N__51605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51594),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52448),
            .ce(),
            .sr(N__51990));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_24_22_6  (
            .in0(N__51567),
            .in1(N__51528),
            .in2(_gnd_net_),
            .in3(N__51516),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52448),
            .ce(),
            .sr(N__51990));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_7 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_24_22_7  (
            .in0(N__52947),
            .in1(N__52941),
            .in2(N__52899),
            .in3(N__52692),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52448),
            .ce(),
            .sr(N__51990));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_0 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_24_23_0  (
            .in0(N__52650),
            .in1(N__52691),
            .in2(N__52869),
            .in3(N__52587),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52441),
            .ce(),
            .sr(N__51994));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_3 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_3  (
            .in0(N__52688),
            .in1(N__52647),
            .in2(N__52588),
            .in3(N__52827),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52441),
            .ce(),
            .sr(N__51994));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_4 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_24_23_4  (
            .in0(N__52646),
            .in1(N__52687),
            .in2(N__52782),
            .in3(N__52586),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52441),
            .ce(),
            .sr(N__51994));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_5 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_5  (
            .in0(N__52690),
            .in1(N__52649),
            .in2(N__52590),
            .in3(N__52731),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52441),
            .ce(),
            .sr(N__51994));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_23_7 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_24_23_7  (
            .in0(N__52689),
            .in1(N__52648),
            .in2(N__52589),
            .in3(N__52536),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52441),
            .ce(),
            .sr(N__51994));
endmodule // MAIN
